Jag måste gå och sova.
Muiriel är 20 nu.
Lösenordet är "Muiriel".
Jag kommer tillbaka snart.
Jag vet inte vad jag ska säga.
Det här kommer aldrig att ta slut.
Du är i bättre form än jag.
Du är i vägen.
Jag tjänar 100 euro om dagen.
Det är för att du inte vill vara ensam.
Jag saknar dig.
Du borde sova.
Det förvånar mig inte.
Av någon anledning så känner jag mig mer levande på natten.
Jag ska skjuta honom.
Varför frågar du?
Jag hittade en lösning, men jag hittade den så fort att det inte kan vara den rätta.
Jag spelar Sudoku då istället för att fortsätta störa dig.
Jag älskar dig.
Jag tycker inte om dig längre.
Alla vill träffa dig. Du är känd!
Jag pratar inte japanska.
Jag kan inte japanska.
Jag talar inte japanska.
Jag ville bara kolla min mail.
Jag ville bara kolla min mejl.
Är det mig du menar?
"Vem är det?" "Det är din mor."
"Lita på mig", sade han.
"Hon gillar musik." "Det gör jag med."
Lektionen börjar inte förrän halv nio.
"Har inte vi träffas någon gång?" frågade eleven.
Skytten dödade hjorten.
Bågskytten dödade hjorten.
Om du inte äter dör du.
"Varför ska du inte åka?" "För att jag inte vill."
Natten är ju ganska lång, eller hur?
Saknade du mig?
Har du saknat mig?
Tack så mycket!
De säger att kärleken är blind.
Matematik är som kärlek – ett enkelt koncept, men det kan bli komplicerat.
Hur lång tid tar det till stationen?
Talar du italienska?
Jag skulle aldrig ha gissat det.
Det skulle jag aldrig ha gissat.
Skulle jag kunna få tala med fröken Brown?
Vad vill du?
Vi uppfattar inte saker som dom är, utan som vi är.
Vi ser inte saker som de är, utan som vi är.
Vi ser inte saker som de är, utan som vi är.
Du ser dum ut.
Jag tror jag ska gå och lägga mig.
Jag heter Jack.
Hur säger du det på italienska?
Jag måste gå och handla. Jag är tillbaka om en timme.
Tack, det var allt.
Skulle du vilja dansa med mig?
Jag skulle vilja stanna en natt.
Öppna munnen!
Är det illa?
Jag har tappat min plånbok.
Jag har tappat bort min plånbok.
"Skicka mig saltet, tack." "Varsågod."
Det är för mycket att göra.
Titta på mig när jag pratar med dig!
Vem vill ha lite varm choklad?
Jag har huvudvärk.
Jag har ont i huvudet.
Ring polisen!
God jul!
Frågan är inte vad jag kan vinna utan vad jag har att förlora.
Jag har så mycket arbete så jag stannar en timme till.
Jag är gift och har två barn.
Vinden avtog.
Jag förstår inte tyska.
Jag ger dig mitt ord.
Jag lovar.
Han är redan en man.
Det är kallt.
Jag är törstig.
Livet är vackert.
Han vill inte att du berättar för honom om ditt sexliv.
Han vill inte att du berättar för honom om ert sexliv.
Han vill inte att ni berättar för honom om ert sexliv.
Han du någonsin ätit en bananpaj?
Hjärnan är bara en komplex maskin.
Den här pingvinungen är så söt!
Det är dags att inse att det är omöjligt. Vi kommer aldrig att klara det.
Allt som är för dumt för att sägas sjungs.
Jag vill inte gå till skolan.
Det regnar.
För sent.
Jag läser boken, medan jag äter.
Hon vill inte prata om det.
Stäng dörren när du går.
Om det inte finns någon lösning, så finns det inte heller något problem.
Finns det ingen lösning, finns det inget problem.
Jag kommer inte att förlora.
För ett ögonblick trodde jag att han hade blivit galen.
Jag vill ha en massage. Jag behöver slappna av.
Det här stället har en mystisk atmosfär.
Hon hade på sig en svart hatt.
Jag vill vara mera självständig.
Jag vill vara mer självständig.
Ja! Jag vann två gånger i rad.
Livet i fängelse är värre än ett djurs liv.
Livet i fängelse är värre än ett djurliv.
Jag skapade en genväg på skrivbordet.
Var är du?
Var är ni?
Jag älskar att resa.
Det är inte viktigt.
Jag bryr mig inte.
Femtiotvå procent av brittiska kvinnor föredrar choklad framför sex.
Coles axiom: Summan av intelligensen på planeten är en konstant; befolkningen växer.
I mörkret är alla katter grå.
Jag vill inte ha den längre.
Hon skulle gärna kommit men hon var på semester.
De bråkade.
Jag åt kaviar.
Gav du dricks?
Glöm inte biljetten.
Hur gick din intervju?
Hur gick det på din intervju?
Jag tror inte mina ögon.
Du har köpt fler frimärken än vad som är nödvändigt.
Du borde inte titta ner på honom.
Ni borde fråga honom om råd.
Du borde fråga honom om råd.
Kan du simma lika snabbt som honom?
Vet du inte att han gick bort för två år sedan?
Vem väntar du på?
Jag tycker att du borde vila; du ser sjuk ut.
Vad vill du göra i framtiden?
Du har friheten att använda detta rum hur du än vill.
Du står näst på tur för en befordran.
Du borde gå till tandläkaren.
Du kom inte till skolan i går.
Du ser blek ut idag.
Du behöver inte ta av dig skorna.
Du ser blek ut.
Du har inte den rätta pondusen som chef för avdelningen.
Vad ska du ha?
Kan du inte tala engelska?
Vad ska du med pengarna till?
Hur länge tänker du stanna här?
Du då?
Vad gör du?
Du är lyckligt lottad som har sådana vänner.
Köpte du den på svarta marknaden?
Är du för eller emot planen?
Du måste bli kvitt den där ovanan.
Du måste göra dig av med den där ovanan.
Du vänjer dig snart vid din nya skola.
Du har druckit tre koppar kaffe.
Ni har druckit tre koppar kaffe.
Du klagar alltid.
Dina föräldrar kom inte, eller hur?
Meg ringde efter dig medan du var borta.
Jag tror inte att din teori håller.
Ditt rum är dubbelt så stort som mitt.
Ditt problem liknar mitt.
Berätta om ditt dagliga liv.
Ditt motiv var beundransvärt, men inte ditt agerande.
Du kan komma och se mig närhelst det passar dig.
Ditt förslag är lite extremt.
Jag är säker på att du lyckas.
Jag behöver inte din hjälp.
Din fråga hör inte till ämnet.
Jag glömde ditt paraply på bussen.
Dina synpunkter är inte av någon vikt alls.
Gör ditt val.
Jag kan inte förstå alls vad det är du säger.
Dina skor är här.
Era skor är här.
Var är din skola?
Var ligger din skola?
Var ligger er skola?
Ditt hus är tre gånger så stort än mitt.
Jag tycker att din engelska har blivit mycket bättre.
Jag tror på dig.
Är din lägenhet väl underhållen?
Du ska få en fin present.
Jag ska göra din nya dräkt.
Jag ser fram emot att träffa dig.
Jag vill att du ska jobba hårdare.
Du äcklar mig.
Han, så som du, är en bra golfspelare.
Vem är din lärare?
Jag hade varit på sjukhuset innan du kom.
Jag behöver dig.
Jag behöver er.
Antingen har du eller han fel.
Dina framgångar beror på dina ansträngningar.
Vem tog hand om hunden medan du var borta?
Vem tog hand om hunden medan ni var borta?
Jag kan inte tacka dig nog för det du gjorde för mig.
Jag hoppas att du aldrig blir kommunist.
Jag stannade hemma i går kväll för att kunna ta emot ditt samtal.
Stunden kommer att komma då du känner dig skyldig för det.
Du förstår inte.
Ni förstår inte.
Kastanjer måste kokas i minst femton minuter.
Jag var hungrig.
Vi kan inte leva utan luft.
Vi kan se tusentals stjärnor på himlen.
Det finns inte ett enda moln på himlen.
Kontrasten mellan himlen och berget är slående.
Inget sött utan svett.
Är Ginza Japans livligaste gata?
Banken tar hand om pengar åt folk.
Varje fredagskväll gick de och drack sig fulla.
Finns det något bord för två ledigt på fredag?
Golden Gate-bron är gjord av järn.
Pengar är roten till allt ont.
Om jag blir rik så kommer jag att köpa den.
Jag är pank.
Ta fram din plånbok.
Guld är tyngre än silver.
Jag har inga pengar på mig.
Guldpriset ändras dagligen.
Finns det några biografer här i närheten?
Hennes ögon blir runda av förvåning.
Till min förvåning så hade han en vacker röst.
En spegel reflekterar ljus.
Är du galen?
Läraren kräver utmärkt gjorda arbeten från hans elever.
Lärare måste förstå barn.
Läraren var tvungen att utvärdera alla elever.
Har du varit i Kyoto?
Fisk, tack.
Och till råga på allt fick jag sparken.
Jag gick en konstkurs i fjol.
Jag odlade tomater förra året och de smakade väldigt gott.
Jag odlade tomater förra året och de var väldigt goda.
Vi gör mjölk till ost och smör.
Vi gör ost och smör av mjölk.
Nöden är uppfinningarnas moder.
En olycka kommer sällan ensam.
Stormen utbrast.
Kom igen! Vi kommer bli sena.
Skynda dig, annars missar du tåget.
Tom skynda dig.
Byggnaden uppe på kullen är vår skola.
Jag är uppe och står igen när mitt ben har läkt.
Rökare sjukskriver sig dubbelt så mycket än vad icke-rökare gör.
Dags att stiga upp.
Studerar du kemi?
Pluggar du kemi?
Din dotter går på droger.
Skulle du kunna säga mig vilken station som ligger närmast ditt arbete är du snäll.
Reglerna kräver att vi alla är närvarande.
Du måste ha tålamod.
Ni måste ha tålamod.
Jag svimmade.
Är du galen?
Tycker du om det?
Glöm det.
Jag träffade ingen på vägen hem.
Vid hemkomsten upptäckte jag inbrottet.
Jag vill inte tillbaka.
Du borde se den här filmen om du får chansen.
Det ligger en sax på bordet.
Konstiga saker hände på hennes födelsedag.
Konstiga saker skedde på hennes födelsedag.
Jag hjälper dig gärna.
Han ser blek ut.
Tvätta ditt ansikte.
Tvätta dig.
Du är röd i ansiktet.
Förespråkare av ökade importavgifter är oense med varandra.
Lätt gånget lätt förgånget.
Du ska inte tro att det kommer att bli enkelt.
Jag minskar på godisätandet.
Jag håller på att dra ner på sötsaker.
Vi lagrade höet i stallet.
Det kalla vädret fortsatte i tre veckor.
Jag fryser. Kan jag stänga fönstret?
Hämta mig en torr handduk.
Lätt gånget lätt förgånget.
Ha det så roligt.
Jag hoppas du har kul.
Jag lärde känna honom när jag var student.
Ingen ut av eleverna var försenade till skolan.
Alla eleverna kommer från USA.
Eleverna har tillgång till dessa datorer.
Två tredjedelar av eleverna kom till mötet.
Eleverna såg alla fram emot sommarlovet.
En student vill träffa dig.
Tre studenter. Här är min studentlegitimation.
Skolan är på gångavstånd från mitt hus.
Skolbarn har förkylningar dubbelt så ofta än vuxna.
Jag tappade bort min väska på väg till skolan.
Dags att gå till skolan.
Det är dags att gå till skolan.
Du hinner inte i tid till skolan.
Människan som slutar lära sig är så gott som död.
Minns du det?
Det råder ingen tvekan om att hon älskar honom, men hon vill inte gifta sig med honom.
Kärnvapen är ett hot mot hela mänskligheten.
Jag vill se gatorna.
Generellt sett lever kvinnor längre än män.
Det haglar i regel om sommaren.
Har du någon hostmedicin?
Har ni någon hostmedicin?
Det är ingalunda lätt att bemästra ett främmande språk.
Var snäll och gå till kirurgavdelningen.
Jag behöver en askkopp.
Företaget kämpar för sin överlevnad.
Vi insisiterar på att det skall hållas ett möte så snart som möjligt.
Mötet sköts upp tills nästa fredag.
Konferensen kommer att hållas i Tokyo.
Mötet varade till 5.
När registrerade de medlemmarnas namn?
Mötet avslutades vid lunchtid.
Vi letar efter en nedgrävd skatt.
Vi måste respektera lokala seder.
Vi döpte min son efter min farfar.
Vi döpte min son efter min morfar.
Vi är benägna att slösa tid.
Vi måste följa spelets regler.
Vi är inte i fara nu.
Vi turades om att köra.
Vi känner till legenden om Robin Hood.
Vi misslyckas att förstå ordets mening.
Vi sprang hela vägen till stationen.
Våra eftersträvningar slutade inte med lycka.
Vår lön är liten, fast vi klarar oss.
Det är inte nödvändigt för oss att närvara vid mötet.
Jag hoppas att vädret klarnar upp innan vi ger oss av.
Jag heter Hopkins.
Jag fick en massa myggbett.
Jag skulle vilja lägga undan mina ägodelar.
Skicka ditt bagage i förväg.
Hanako har glömt sitt paraply igen.
Mars är desto mer intressant för dess närliggande likhet med vår jord.
När elden brast ut sov han död som en sten.
Eld är väldigt farligt.
Känner du till kabuki?
Låt oss sjunga och dansa.
Jag är ledig.
Jag orkar inte lyssna mer på hennes klagomål.
Det tog dem två år att bygga huset.
Huset brann ner till grunden.
Jag har spenderat mycket pengar på mitt hus.
Huset brinner.
Tycker du om sommaren?
Tycker du om sommar?
Sommaren är över.
Vem tror du att du är?
Han betonade att tiotusentals människor skulle komma till konserten.
Hur många ingenjörer deltog i konferensen?
När kommer du att vara tillbaka?
Vad läser du?
Så blå himlen är!
Kommer du att lyckas med att reparera min bil?
Vi diskuterade vad vi skulle göra.
Jag vill dricka något kallt.
Har du gjort något nyårslöfte?
Snälla ge mig någonting att äta.
Ge mig något att skriva på.
Kan jag hjälpa dig?
Kan jag hjälpa dig?
Vad vill du att jag ska göra?
Vad är orsaken?
Oavsett vad som händer kommer jag aldrig att ändra mig.
Hur är läget?
Vad händer?
Vad är det som saknas?
Vad saknas?
Vad är det där borta?
Vad fick dig att komma hit?
Håll mig informerad tack.
Få saker ger oss så mycket nöje som musik.
Hade jag fel?
Det finns ingenting jag kan göra.
Jag pratar inte med dig; jag pratar med apan.
Lämna mig ifred!
Låt mig vara!
Det är min CD-skiva.
Det är min CD.
Titta på huset med det röda taket.
Jag såg månen ovanför taket.
Länge leve konungen!
I Europa och Amerika ser de hunden som en familjemedlem.
Sluta göra omsvep och kom till saken.
Sluta gå som katten kring en het gröt och kom till saken.
Segla längst kusten.
Jag växlade yen till dollar.
Det är en timmes promenad till stationen.
Stationen är två engelska mil bort.
Finns det en bank nära stationen?
Finns det någon bank nära stationen?
Kan du hämta mig på stationen?
Kan ni hämta mig på stationen?
Väntar du på oss vid stationen?
Väntar du på oss på stationen?
Väntar ni på oss på stationen?
Väntar ni på oss vid stationen?
Kommer du att vänta på oss på stationen?
Kommer du att vänta på oss vid stationen?
Kommer ni att vänta på oss vid stationen?
Kommer ni att vänta på oss på stationen?
Var inte rädd för att göra misstag när ni pratar engelska.
Låt oss tala engelska.
Engelska är svårt, inte sant?
Engelska är svårt, eller hur?
Engelska talas i många länder runt om i världen.
Engelska är, som du vet, i högsta grad ett levande språk.
Engelska är, som ni vet, i högsta grad ett levande språk.
Hur många engelska ord kan du?
Att simma över sjön tog nästan kol på mig.
Jag var på bio.
Filmen börjar klockan tio.
Filmen var intressant, precis som jag hade förväntat mig.
Föraren svängde ratten till höger.
Det har slutat att regna.
Det har slutat regna.
Regniga dagar gör mig deppig.
Trots att det regnade ställdes matchen inte in.
Regnet slog emot fönstren.
Jag kanske går ut om det slutar regna.
Regnet föll i mitt ansikte.
När det slutar regna ska vi ta en promenad.
Jag kan inte böja min högerarm.
Jag kan inte se något med mitt högra öga.
Ligg på din högra sida.
Jag har en ärta i min högra näsborre.
Din högra strumpa är utochinvänd.
Ett högt träd kastar sin långa skugga på vattnet.
Å ena sidan är han snäll men å andra sidan är han lat.
För Amerikaner, på andra sidan, är det mer troligt att ta risker i hopp om att uppnå stora framgångar.
Vad i hela världen står på?
Om han ansträngde sig så skulle han lyckas.
Jag tänker så det knakar, men jag kan inte komma på hennes namn.
Jag ogillar att vara ensam.
En man kom fram till mig och bad om en tändsticka.
Låt mig vara.
Lämna mig ifred.
Vill du följa med?
Jag gillar inte att bli driven med.
I medicinsk forskning är en av de största problemen att isolera orsaken till sjukdomen.
Vad sa han?
En sexsiffrig inkomst är inte ovanligt för en läkare.
Jag fick en bot på tjugo dollar för olovlig parkering.
Min mage kurrar.
Jag förlorade medvetandet.
Kommittén sammanträder två gånger om månaden.
Kommittén sammanträder två gånger i månaden.
Kommittén sammanträder två gånger per månad.
Jag brukade inte röka.
Det brukade finnas en restaurang framför den här busstationen.
När man talar om trollen står de i farstun.
Han är helt hopplöst dålig.
Det jag inte vill förlora är kärlek.
Vi måste försöka bryta dödläget.
Jag måste göra klart läxan innan middagen.
Jag föredrar att åka tåg framför att flyga.
Jag vill gå med dig.
Jag är från Kyoto.
Jag är så lycklig!
Jag hann dit i tid.
Jag har en vän vars far är en känd pianist.
Verkligen. What kan jag göra?
Klockan är sju i London nu.
Hon är sju i London nu.
Långa kjolar är på modet.
Rock tilltalar unga män och kvinnor.
Vi skulle vilja ha en flaska rosé.
Raketen är i omloppsbana runt månen.
Håll i repet.
Håll repet.
Kan du släcka ljusen?
Kan du släcka stearinljusen?
Roy behövde inte skynda sig till flygplatsen för att möta hans föräldrar.
Kan jag köpa enbart linserna?
När måste jag lämna in rapporten?
Lucy kan inte använda ätpinnar.
Lucy är en fin liten flicka.
Lynn springer snabbt.
Linda älskar choklad.
Jag skulle vilja ha två kilo äpplen.
Snälla ta det lugnt.
Snälla lugna ner dig.
Vilken tid avgår bussen till flygplatsen?
En bra lärare måste vara tålmodig med hans elever.
En ekorre gömde sig bland grenarna.
Lejonet öppnade sin enorma mun och vrålade.
Lejonet är kungen av djungeln.
Jag ser honom ofta.
Jag träffar honom ofta.
I Europa startar skolorna i september.
Låt oss hoppas på bra resultat.
Ha en bra dag.
Ta din tid.
Jag var missnöjd över att det fanns så lite att göra.
Bergets övre del är snötäckt.
Det kanske blir regn snart.
Kärleken kommer så småningomg
Prata långsammare.
Ät mer, annars kommer du inte att få styrka.
Jag önskar att vi hade mer tid.
Du borde äta mer frukt.
Vill du ha mer kakor?
Vad skulle du göra om du såg ett spöke?
Vad skulle hända om han skulle komma försent?
Om det regnar kommer han inte.
Om jag visste hennes namn och adress kunde jag skriva till henne.
Om ni har något problem så fråga mig om hjälp.
Om jag vore en fågel så skulle jag kunna flyga till dig.
Har du inga pengar så får du klara dig utan.
Jag gör det om du stöttar mig.
Jag ber om ursäkt om jag har sårat dig.
Jag är så mätt.
Du kan lämna rummet nu.
Har du ringt henne än?
Det är dags att du börjar stå på dina två egna fötter.
Har du ätit lunch än?
Snälla sänk volymen lite till.
Vill du ha lite mer nötkött?
Våren är kommen.
Jag måste gå nu.
Jag måste bege mig nu.
Jag måste bege mig nu.
Jag måste bege mig nu.
Vi ska ha barn.
Jag kan inte vänta längre.
Det är bäst att du inte väntar längre.
Har far kommit hem ännu?
Det är dags för mig att gå.
Kan du säga det en gång till?
Försök igen.
Mary och Jane är kusiner.
Det har blivit märkbart kallare.
Meg köpte en burk tomater.
Meg pratar för mycket.
De talar spanska i Mexiko.
Mary ser ovänlig ut, men egentligen har hon ett gott hjärta.
Mary sprang.
Hur mår Mary?
Mary kan simma.
Mary gillar mjölk väldigt mycket.
Mary är en väldigt söt tjej.
Mary har all anledning att vara nöjd.
Alla hoppades att hon skulle vinna.
Jag mindes alla.
Tala högre så att alla kan höra dig.
Mjölken kokade över.
Mjölken surnade.
Kortkorta kjolar har blivit omoderna.
Damer och herrar, välkomna ombord.
Hon ser ut att vara full.
Mayuko kan cykla.
Mayuko verkar klok.
Det tog inte lång tid innan månen kom fram.
Jag skrev till honom av en helt annan anledning.
Jag har fortfarande inte funnit det jag söker efter.
Jag har fortfarande inte hittat det jag letar efter.
Har du inte bestämt dig än?
Låt oss göra det någon annan gång.
Först och främst måste vi bestämma oss för ett namn.
Först och främst måste du leta upp det i ordboken.
Inte så mycket senap.
Moder Teresa föddes 1910 i Jugoslavien.
Du måste skörda det du har sått.
Hur mår du, Mike?
Jösses, vilken oanständig kund!
Herr White är en förnuftets man.
Herr White är en förnuftig man.
Här är hon!
Här kommer han.
Bob har många böcker på sitt rum.
Har Bob rätt?
Bob är min vän.
Bob är min kompis.
Bob var inte med på planen.
Bob tittade förbi hos sin farbror.
Vi börjar mötet när Bob kommer.
I de flesta fall likställs modernisering med västernisering.
Finns det något vatten i kannan?
En av dina knappar har lossnat.
Se upp för ficktjuvar.
Jag vill ha lite pengar.
För egen del föredrar jag kaffe framför te.
Själv föredrar jag kaffe framför te.
Jag har inte råd att betala så mycket.
Var är de andra flickorna?
Vill du beställa någonting mer?
Var någon annan frånvarande?
Vem mer kom till festen?
Tror du vi hinner i tid till flygplatsen, Paul?
Paula måste hjälpa hennes pappa i köket.
Ben har också något med saken att göra.
Han satte sig på bänken.
Vi blev stupfulla.
Helen håller alltid sitt rum rent.
En helicopter åkte runt över oss.
Vem har vi att tacka för penicillinets upptäckt?
Betty gick till havet i går.
Min katt dog igår.
Bess är endast ett barn.
Ge mig en flaska vin.
Det saknas en gaffel.
Vad är Finlands huvudstad?
Bill hatar att hans far röker mycket.
Bill lyckades bli godkänd på provet.
Bill är på väg till New York.
Bill, ring mig ikväll.
Det ser ut som att det ska börja regna.
Det ser ut att bli regn.
Den ena talar engelska, den andra japanska.
Det fanns inte en själ i sikte.
Jag har en idé.
Jag hade en besvärlig tid.
Jag hade det besvärligt.
Det var ett förskräckligt väder.
Jag har slutat med öl.
Peter är inte alls lik hans pappa.
Peter ser väldigt ung ut.
Ett piano är dyrt.
Bröd bakas i ugn.
Bröd bakas i en ugn.
Hawaii har fint väder året runt.
Låt oss spela volleyboll.
Det är femtio kilometer till Paris.
Jag funderar på att åka till Paris.
Var ligger Paris?
Harry är bara 40.
Patricia kommer att hålla i turneringen.
Ingen väntar vid busshållplatsen. Vi kanske har missat bussen.
Jag går hellre än att ta bussen.
Någon stal mitt pass.
Vi hade det väldigt svårt att hitta busshållplatsen.
Vi hade stora svårigheter att hitta busshållplatsen.
Ta en buss.
Hur kan jag åka buss till sjukhuset?
Byron lämnade England för att aldrig komma tillbaks igen.
Jag letar efter ett deltidsjobb.
Vi välkomnar alla som vill komma till festen.
I länder som Norge och Finland har de mycket snö på vintern.
Har du någonsin hört talas om Nessie?
Råttor förökar sig fort.
En fladdermus är lika lite fågel som en råtta.
Morötter och rovor är ätbara rötter.
Staten New York är nästan lika stort som Grekland.
Hur stor är New York Citys befolkning?
New Yorks gator är väldigt breda.
Vad?
Vilken spännande match!
Åh nej! Mitt hus brinner!
Vilken vacker fågel det är!
Vad vill du att jag ska prata om?
Nancy handlade lite på vägen.
Nancy tycker om inomhussporter.
Visst är han ung, men han är mycket pålitlig.
Han må vara ung, men han är verkligen en tillförlitlig person.
Det stämmer att projektet är en svår uppgift, men herr Hara kommer att kunna göra det.
Varför är du arg på honom?
Varför kommer du så tidigt?
Varför uppför sig män som apor, och vice versa?
Varför ser du så ledsen ut?
Varför?
Varför är du så trött idag?
Vi måste kompensera för den förlorade tiden.
Jag kunde inte somna.
Vad gör den här stolen här?
Ah, föraren är galen.
Ingen medicin kan bota denna sjukdom.
Ingen medicin kan bota den här sjukdomen.
För vilken anledning bröt du dig in i huset?
Vilken sorts vin rekommenderar du?
Vilken typ av sport gillar du?
Varje moln har en silverkant.
Vilken säng som helst är bättre än ingen säng alls.
Oavsett hur snabbt du kör hinner du inte dit i tid.
Tom slog ner honom.
Tom är inte en lat pojke. I själva verket arbetar han hårt.
Tom är inte här.
Tom är frånvarande.
Tom ser blek ut.
Tom arbetade hårt bara för att misslyckas på tentan.
Var är Tom född?
Tom förlöjlar sig alltid över John på grund ut av hans dialekt.
Tom gör alltid narr ut av John på grund ut av hans dialekt.
Tom hittar alltid fel hos henne.
Var är Toms klassrum?
Tom har många talanger.
Tom är förlovad med Ruth.
Är inte du Tom?
Stör inte Tom medan han läser.
Jag ska prata med Tom när han kommer hem.
Vem vikarierar för Tom medan han är borta?
Vilken tunnelbanelinje går till stadskärnan?
Vilken tunnelbanelinje går till centrum?
Alla sittplatser var upptagna.
Vilken ordbok syftade du på?
Var gör det ont?
Vilken frukt tycker du bäst om?
Hur lärde du känna henne?
Du kan alltid räkna med honom i ett nödfall.
Hur länge har du varit utomlands?
Vad kostar det?
Hur långt kommer det att ta för att bli återställd?
Vilken bra tennisspelare Tony är!
Var är Tony?
Det var väldigt svårt.
Det är skönt och varmt.
Trots kylan gick vi ut.
Jag känner mig väldigt kall.
Vilket som. Det är oviktigt.
Vem vinner?
Vart skulle du vilja åka?
Du kan välja vilken bok du vill.
Ni får välja vilken bok som helst.
Det spelar ingen roll vilket lag som vinner matchen.
Vem arbetar du för?
Du kan välja vilken du vill.
Vilken är din gitarr?
Förresten, hur många av er för dagbok?
Förresten, spelar du fiol?
Förresten, var bor du?
Var bor du, förresten?
Hur gammal är du egentligen?
Var får jag tag på böcker?
Var arbetar du?
Var kan jag köpa frimärken?
Var ska vi träffas?
Var ska vi ses?
Det är en bra regel varsomhelst att se åt båda håll innan du gå över gatan .
Mår du inte bra?
Jag undrar vem som satte igång det där ryktet.
Kan du komma?
Förlåt.
Jag fattar inte.
Varsågod och ta lite tårta.
Varför kommer hon inte?
Vad hände? Bilen saktar ner.
Vad fattas dig? Du ser blek ut.
Kan jag få ett glas vatten, tack.
Jag kan inte prata tyska.
Tyskan är inte ett lätt språk.
Stäng dörren.
Dörrar är inte så illa som du tror.
Pojken som står vid dörren är min bror.
Kan du vara snäll och låsa dörren?
Kan ni vara snälla och låsa dörren?
Kan du låsa dörren är du snäll?
Kan ni låsa dörren är ni snälla?
Jag hörde dörren stängas.
Var snäll och stäng av teven.
Mary gillar att titta på TV.
Skruva ner tv:n.
Tack vare televisionen är pojkar och flickor benägna att ej läsa böcker.
Jag såg en gammal film på tv.
Jag tror inte att tv någonsin kommer att ersätta böcker.
Men det var förstås länge sedan.
Jag spelar en timmes tennis varje dag.
Jag spelar tennis en timme om dagen.
Dennis kan göra det fulaste grimasen i staden.
Jag är säker på att Teds hostande beror på rökning.
Kom ner så snart som möjligt.
Jag lämnar tillbaka boken så fort jag kan.
Texas är nästan dubbelt så stort som Japan.
Katten på bordet sover.
Det ligger en bok på bordet.
Jag kanske har lagt den på bordet.
Det finns ett äpple på bordet.
Jag hittar inte Tim.
Äter du ofta fisk till middag?
En efter en reste sig och gick.
Jag kollade på klockan och visste vilken tid det var.
Var snäll och vänta en stund medan jag gör klart ditt kvitto.
Ge mig tre kritor.
Jag ska strax gå.
Jag är inte det minsta orolig.
Kyckling, tack.
Jag ska lära dig att spela schack.
Jag vill köpa en tjeckisk tröja.
Dagarna blir längre och längre.
Dagarna blir allt längre.
Tankfartyget har bara en liten besättning ombord.
Ingen sprang före honom.
Ingen kan lyckas med något utan ansträngning.
Vem som helst kan göra misstag.
Alla verkar gilla golf.
Vi behöver alla acceptera flödet i dessa tider.
Det är ingen tvekan om vem som blir vald.
Vem har skrivit denna bok?
Kan någon öppna den här dörren, tack?
Det luktar som om någon har rökt här inne.
Någon verkar ropa på mig.
Någon måste ha tagit mitt paraply av misstag.
Hon kommer förmodligen.
Han kan mycket väl ha rätt.
Han kan ha rätt.
Det kommer att regna.
Han har kanske många flickvänner.
Varför slutar du inte röka?
Du får inte röka.
Ni får inte röka.
Hon målar varje dag, oavsett hur mycket hon har att göra.
Det tog nätt och jämnt en timme.
Skulle du kunna förklara vägen till Madame Tussaud?
Skulle ni kunna förklara vägen till Madame Tussaud?
Han har gått till Nagoya för affärer.
Att flyga drake kan vara farligt.
Många människor dödades i kriget.
Dykarna hittade ett skeppsvrak på havsbottnen.
Låt oss inte tänka så.
Du får inte beté dig så.
Det är dumt att läsa en sådan tidskrift.
Det där är en bit paj.
Det är bara en ursäkt.
Det är onormalt att äta så mycket.
Jag uppfattade inte riktigt namnet på den där designern.
Jag ger mig av nu.
Det är dags att börja röra mig härifrån.
Stäng av den.
Man har inte hört något ifrån dom sen dess.
Har du varit här sen dess?
Varför letar du inte upp det i telefonkatalogen?
Kan du bevisa det?
Låt mig se det där.
De är min farfars böcker.
De är min morfars böcker.
Vad är de gjorda av?
Det är ungefär lika stort som ett ägg.
Det är en sjukdom som inte kan förebyggas.
Det kan inte vara sant.
Det visade sig vara sant.
För henne är det en förolämpning.
Det var ett misstag från deras sida.
Det kommer att kosta minst fem dollar.
Det är en bild som jag gillar väldigt mycket.
Betyder det att du vill göra slut?
Jag kanske gör det; det beror på omständigheterna för tillfället.
Det är enkelt att göra och det är billigt.
Det är bara ett talesätt.
Det är upp till dig.
Oj! Det är billigt!
Det är värt ett försök.
Det var ett väldigt spännande spel.
Det är ett för svårt problem för mig att lösa.
Det är skräp. Släng det!
När börjar det?
Vad menar du med "den"?
Jag vet inte vad det är.
En lång tystnad följde.
Jag heter inte "flicka" heller.
Vad betyder det?
Här är bussen.
Gubben är blind på ena ögat.
Den gamle mannen är blind på ena ögat.
Den gamle mannen satte sig ner.
Den gamle mannen var inte så elak som han såg ut att vara.
Den väljaren, Mary Johnson, visade sig vara demokrat.
Medicinen gjorde underverk för hans hälsa.
Medicinen smakar beskt.
Drogens effekter är intensiva men kortvariga.
De goda nyheterna fick henne att gråta.
Jag har läst ut boken.
Lägg tillbaks boken där du fann den.
Juvelen stals under natten.
Soldaten uppgav sitt namn.
Soldaterna var utrustade med vapen.
Ljudet väckte mig från min sömn.
Ljudet kommer att väcka bebisen.
Ingen kunde förklara hur saken var gjord.
Fången var bakom galler i två månader.
Varför provade du inte klänningen innan du köpte den?
Satte du på frimärket på brevet?
Rummet är fullt av folk.
Min bror och jag delade rummet.
Jag hittade rummet tomt.
Har rummet ett badkar?
Rummet städas av fru Smith.
Rummet kommer att målas imorgon.
Det fanns ingen i rummet.
Det var en massa möbler i rummet.
Rummet har två fönster.
Det fanns nästan ingenting i rummet.
Det finns ett piano i rummet.
Det finns en TV i rummet.
Det finns två hundra personer i rummet.
Damen förblev tyst.
Damen är över åttio.
Paret hade ett lyckligt liv.
Fastighetsmäklaren ljög för paret.
Fyll flaskan med vatten.
Den stackars mannen blev äntligen en känd artist.
Den sjuka mannens liv är i fara.
Sjukhuset öppnade förra månaden.
Isen är väldigt tjock.
Ord kan inte beskriva skönheten.
Den vackra kvinna är vänlig.
Planet flög över Mt. Fuji.
Planet gjorde en perfekt landning.
Flygplanet lyfte för tio minuter sedan.
Det var femtio passagerare på planet.
Dörren öppnar nu.
Dörren är öppen nu.
Tjejen är ensam.
Jag är säker på att jag rätt nummer.
Det var väldigt kallt den kvällen.
Jag kan inte stå ut med ljudet.
Uppfinnaren är känd över hela världen.
Ta bort lådan.
Titta inte in i lådan.
Lådan är för tung för att lyftas.
Lådan är nästan tom.
Lådan var nästan full.
Det är en massa ägg i lådan.
Lägg ingenting på lådan.
Vad finns i lådan?
Lådan var full av böcker.
Det fanns ingenting i lådan.
Katten klängde vid hennes klänning.
Det var kallt hela den dagen, och senare började det regna.
Svaret är helt fel.
Flygfältet på ön är nu täckt med ogräs.
Jag håller inte med dig på den punkten.
Affären är öppen året runt.
Affären är öppen året om.
Trädgården har blivit proffesionellt anlagd.
Kämpa!
Staden förstördes under kriget.
Skulpturerna är av högt värde.
Koppen är sprucken.
Var kan jag få tag på kartan?
Jordbävningen skakade husen.
Vi har väldigt besvikna över att höra nyheterna.
Killen var så barnslig att han inte kunde motstå frestelsen.
Mannen erkände slutligen vad han hade gjort.
Mannen erkände äntligen vad han hade gjort.
Mannen erkände till slut vad han hade gjort.
Mannen erkände till sist vad han hade gjort.
Pojken tömde tallriken på ett ögonblick.
Virvelvinden tog med sig förlust av regn till det distriktet.
Vi såg båten gungande ute på den stormiga sjön.
Floden är femtio meter vid.
Jag tvättade medan spädbarnet sov.
Spädbarnet döptes till Alfred efter sin farfar.
Spädbarnet döptes till Alfred efter sin morfar.
Båda eleverna klarade av alla prov.
Den nya maskinen kommer att ta upp en massa utrymme.
Sex blev inbjudna, inklusive pojken.
Sex var inbjudna, pojken inkluderad.
Pojken gick vilse i skogen.
Pojken gjorde sig lustig över flickan.
Det var snudd på otänkbart att pojken skulle stjäla.
Flickan stirrade på dockan.
Hyddan stacks i brand.
Kojan stacks i brand.
Skjulet stacks i brand.
Skådespelerskan har ett väldigt vackert namn.
Så fort som tjejen såg sin mamma så började hon att böla.
Flickan gick in i rummet.
Inrättningen måste skyddas.
Vem skrev brevet?
Bilen förbrukar mycket bränsle.
Frågan var omöjlig för oss att besvara.
Inte förrän då fick han reda på sanningen.
Endast då förstod jag vad han menade.
Välgörenhetsorganisationen har fått sitt namn efter en man som donerade cirka 2 miljarder yen.
Ingen kan förneka detta faktum.
Olyckan skedde i det hörnet.
Det tjänar inget till att bråka med honom om det.
Direktören gav exakt det svaret som jag letade efter.
Barnet tigger alltid om någonting.
Det tog henne hela eftermiddagen att göra klart arbetet.
Det är svårt att utföra uppgiften.
Arbetet är nu igång.
Den internationella konferensen skulle gå av stapeln i februari i år.
Landet förklarade krig mot sitt grannland.
En revolution bröt ut i det landet.
Vad betyder det här ordet?
Sjön är stor och vacker.
Isen över ån är för tunn för att kunna bära din vikt.
Det bodde en gubbe i det gamla huset.
Det bodde en gammal man i det gamla huset.
Det bodde en gammal gubbe i det gamla huset.
Hunden är döende.
Hunden grävde en grop.
Hunden vill gå ut.
Hunden är på stolen.
Hunden heter Ken.
Gå inte nära hunden.
Följden blev att hon förlorade jobbet.
Planen stöddes av praktiskt taget alla närvarande.
Festen hölls i professorns ära.
Tåget bör vara i Osaka vid tio.
Skrivbordet är av trä.
Det underliga ljudet fick henne upp ur sin säng.
Skolan ligger en halv mil iväg från mitt hus.
Skolan ser ut som en fängelse.
Den här skolan grundades år 1970.
Klippan är nästan vertikal.
Bilden är verklighetstrogen.
Bilden kostar tio pund.
Nyhetsförmedlaren betonar matkrisen för mycket.
Företaget vill anställa 20 personer.
Företaget gick i konkurs.
Företaget bidrar med sjukvård och livförsäkringar åt alla dess anställda.
Låten var en stor succé.
Huset höll på att målas av min far.
Huset är målat i vitt.
Huset omgavs av en stenmur.
Musikern är känd i utlandet såväl som i Japan.
Oljuden väckte mig.
Jag tar den gula.
Det var du som föreslog att vi skulle se den filmen.
Doktorn funderar noggrant innan han bestämmer sig för vilken medicin han ska ge.
Hönan har värpt ett ägg.
Hotellet drivs av hans farbror.
Hotellet drivs av hans morbror.
Hotellet har en bra utsikt.
Båten lade till nära kusten.
Sitt inte på den där bänken är du snäll.
Festivalen kommer att gå av stapeln nästa vecka.
Öppna flaskan.
Byggnaden totalförstördes i jordskalvet.
Den slipsen passar dig tillsammans med din skjorta.
Det tar oss fem minuter att gå igenom tunneln.
Det händer att dörren är öppen ibland.
Var köpte du biljetten?
Diamanten värderades till 5 000 dollar.
Soporna ger ifrån sig en förfärlig stank.
Tappa inte den där koppen.
Kaffet var så varmt så jag inte kunde dricka det.
Det är roligt att spela baseball.
Gruppen springer på stranden.
Vi såg inga flickor i gruppen.
Spiken gick igenom väggen.
Kragen sitter åt för hårt runt min hals.
Jag ångrar att jag åt ostronen.
Hissen verkar vara trasig.
En del av uppsatserna är mycket intressanta.
Jämför de båda noggrant, så ska du se skillnaden.
Jag åkte dit med buss och tåg.
Där är Tokyo.
Det var ingen där förutom jag.
Det fanns ingen där förutom jag.
Det tar inte särskilt lång tid.
Jag är inte trött alls.
Jag är inte ett dugg trött.
Jag är inte alls trött.
Denna stol är ful.
Den här stolen är ful.
Du borde ha besökt Kyoto.
Ursäkta, kan du förklara vägen till stationen?
Skulle du kunna sänka radion?
Herr Smith gläder sig över sin sons framgång.
Herr Smith har gjort det till en regel att ta en promenad varje morgon.
Det beror helt på huruvida de kommer att hjälpa oss.
Alla människor andas luft.
Alla pojkarna sprang iväg.
Jag är nöjd med allt.
Jag får svår prestationsångest före jag ska hålla ett tal.
Jag har redan sagt det till dig.
Jag kommer.
Jag kommer tillbaka snart.
Genast lämnade fåglarna sina bon.
Du kan lika gärna börja omedelbart.
Du kan lika gjärna lämna hemmet på en gång.
Jag kan åka skidor.
Sveriges befolkning ökar.
Sverige har sitt eget språk.
Schweiz är beläget mellan Frankrike, Italien, Österrike och Tyskland.
John byggde en bokhylla.
John borde vara här när som helst nu.
John er mun hærri en Mary.
John är bra på schack.
John gillar schack.
Jag tycker om schack.
John kan inte göra det, och inte jag heller, och inte du heller.
John sitter vid Jack.
John sitter bredvid Jack.
John spelade gitarr och hans vänner sjöng.
John är här om fem minuter.
John's mor ser så ung ut så att hon ofta misstas för en ut av hans äldre systrar.
Jo-Jo var en man som trodde att han var en ensamvarg.
Jag letar efter något att tvätta mattan med.
Sen då?
Jag kan inte stänga av duschen. Kan du kolla det åt mig?
Jag lyckas inte stänga duschen. Kan du kolla på det åt mig?
Jag måste stryka min skjorta.
Jack samlar på frimärken.
Jack kan engelska.
Jack då?
Det var fönstret som Jack tog sönder igår.
Jim kommer inte bra överens med sina klasskamrater.
Jimmy insisterade på att jag skulle ta honom till zoot.
Låt mig fundera ett litet tag.
Gå in och vinn!
Men hon tyckte om barn och gillade sitt jobb.
Men snart skulle han inte kunna gå, skriva eller ens äta själv.
Men han ville väldigt gärna ha en son.
Jane ska undervisa våra elever från och med nästa vecka.
Jane är fet, ohövlig och röker för mycket. Men Ken tycker att hon är förtjusande och härlig. Det är därför de säger att kärleken är blind.
Det är möjligt att Jane inte är hemma just nu.
Vad gjorde Jean?
Har Jane lämnat Japan för gott?
Jane spelade väl inte tennis?
Det här halsbandet som tillhör Jane är en gåva från hennes mormor.
Det här halsbandet som tillhör Jane är en gåva från hennes farmor.
Ingen dramatiker kan jämföras med Shakespeare.
Fotboll är inte nödvändigtvist begränsat till män.
Fotboll är populärare än tennis.
Du måste vara jättehungrig nu.
Amen ge dig iväg.
Är du redo att beställa nu?
Är ni redo att beställa nu?
Det är fritt för fantasin.
Eftersom varorna Ni debiterat oss inte var perfekta kommer vi inte att betala räkningen.
Tusen tack för din vänlighet.
Tusen tack för er vänlighet.
Jag kommer inte att glömma bort din vänlighet så länge jag lever.
Jag uppskattar verkligen dina råd.
Jag önskar dig ett lycka till.
Jag är tacksam för din hjälp.
Jag är tacksam för er hjälp.
Vill du göra mig sällskap?
Datorn jämförs ofta med människans hjärna.
Du hade inte behövt köpa ett sådant stort hus.
Jag vill komma ut härifrån!
Du borde inte gå ut i den här kylan.
Du kan inte förvänta dig en sådan bra chans igen.
När det regnar såhär får vi aldrig en chans att gå!
Jag trodde aldrig att ett såhär fint hotell skulle finnas på en sådan här plats.
Sydde du den här för hand?
Får jag prova den här?
Vem förstörde denna?
Vem förstörde det här?
Kunde du ta det här, tack?
De här verktygen behövs verkligen repareras.
Kan du visa mig en billigare kamera än denna?
Så här långt ser det bra ut.
Detta är deras hus.
Detta är huset där han bor.
Detta är en kamera tillverkad i Japan.
Det här är den vackraste blomman i trädgården.
Det här är ett sådant enkelt problem så att vilken elev som helst kan lösa det.
Det här är en liten bok.
Det här är en bild av min syster.
Det här är min väska.
Det här är den vackraste utsikten som jag någonsin sett.
Det här är det sötaste spädbarnet jag någonsin har sett.
Detta används fortfarande dagligen.
Det här är ett mycket märkligt brev.
Det här är en mycket märklig bokstav.
Det här är en läsvärd bok.
Det här är en penna.
Kan du förklara vad det här är?
Var det här någon annans idé?
Det är just den boken som jag har väntat så länge på för att läsa.
Det här är just den ordbok jag har letat efter.
Det är just den här ordboken som jag har letat efter.
Jag behöver en låda i den här storleken.
Det här är ett postkontor och det där är en bank.
Det här är det värsta av allt.
Jag är inte säker på om det här är rätt.
Detta är min bil.
Detta är huset jag bodde i när jag var barn.
Här är mitt kvitto.
Bara du kan göra detta.
Det här är roten till problemet.
Är det din bok, Mike?
Gillar du golf?
Förlåt, men jag hör dig ej så bra.
Förlåt, det var inte min mening att sparka dig.
I den här tidningen avgränsar jag diskussionen om Emmets 'dyad' stil i hans verk 1995.
Det här tåget går mellan Tokyo och Hakata.
I hur många minuter ska jag koka den här frusna sparrisen?
Det här ägget är färskt.
Inga av de här äggen är färska.
Posta det här brevet.
Den här medicinen kommer att bota din förkylning.
Det är inte lönt att försöka lösa det här problemet.
Det är ingen mening med att försöka lösa det här problemet.
Vi behöver tänka över problemet mer försiktigt.
Den här boken behandlar Kina.
Den här boken innehåller fyrtio fotografier.
Den här boken är tung.
Den här boken tillhör mig.
Den här boken finns bara tillgänglig i en affär.
Denna bok duger.
Den här boken duger.
Finns det en bank i närheten?
Finns det en bensinmack i närheten?
Den här klänningen skrynklar sig lätt.
Det här rummet är allt annat än varmt.
Det här tyget känns lent.
Håller isen?
Vad finns i den här lådan?
Du måste ta tjuren vid hornen!
Sammanfatta innehållet i 60 engelska ord.
Den här vägen kommer att leda dig till parken.
Följ den här gatan i ungefär fem minuter.
Hur bred är den här vägen?
Den här genomskinliga vätskan innehåller gift.
Denna genomskinliga vätska innehåller gift.
Det har varit en mycket svår vinter.
Denna punkt är värd att betona.
Denna punkt förtjänar särskild emfas.
Vi kan inte hålla med dig på denna punkt.
Den här pojken har en stark, sund kropp.
Jag står inte ut med det här oljudet längre.
Är det säkert att simma i den här floden?
Kan jag avboka den här biljetten?
Den här stenen är dubbelt så tung som den där.
Är den här platsen upptagen?
Denna produkt är tillverkad i Italien.
Den här produkten är tillverkad i Italien.
Det här vattnet smakar bra.
Den här maten luktar ruttet.
Jag vill sända detta paket till Canada.
Den här romanen är översatt från engelska.
Vem är det som äger pistolen?
Olyckor av det här slaget sker ofta.
Den här sortens arbete kräver mycket tålamod.
Den här pjäsen har ingen humor i sig.
Det här gräset behöver klippas.
Den här bilen drivs av alkohol.
Den här bilen går på alkohol.
När kan jag se dig igen?
Jag kompenserar för det nästa gång.
Den här klockan verkar inte fungera som den ska.
Den här tanden sitter löst.
Du kan använda ett lexikon till den här tentamen.
Detta barnet har växt upp normalt.
Jag tror inte att ungen kom till Tokyo själv.
Det här arbetet är inte på något sätt lätt.
Jag tar det här paraplyet.
Du borde rensa ogräset.
Det finns många städer i det här landet.
Den här gamla fisken smakar konstigt
I det här fallet tror jag att han har rätt.
Den här dramaserien kommer att sändas imorgon.
Det kommer att ta några dagar att gå in de här skorna.
De här kängorna tillhör henne.
Dom här skorna är dyra, och dessutom är dom för små.
De här skorna är en aning för stora.
De här skorna sitter inte särskilt bra.
De här skorna är gjorda i Italien.
Dessa skor är tillverkade i Italien.
Det finns inga matbutiker i närheten.
Den här bron byggdes för två är sedan.
Det här klassrummet är städat.
Det här monumentet restes i februari 1985.
Den här maskinen går på elektricitet.
Gå upp för den här trappan.
Den här firman trycker många läroböcker.
Jag skulle vilja skicka dessa till Japan.
De här blommerna blommar tidigare än vad andra gör.
Det är farligt att bada i den här floden.
Den här sången är en kärlekssång.
Den här låten påminner mig alltid om mina skoldagar.
Det här huset behöver målas.
Det här kommer att bli den varmaste sommaren på trettiosex år.
Den här filmen är sevärd.
Den här roboten gör vad jag än säger. Det är till stor hjälp när jag är för trött för att göra någonting. Inte alltför troligt, va?
Vad kostar den här radion?
Sådant kan hända då och då.
Städa golvet med den här moppen, tack.
Mjölken håller i två dagar.
Den här gammla bilen går sönder hela tiden.
Denna salen tar 2000 personer.
Du får inte formatera den här disketten.
Det här vinet smakar gott.
Det här vinet är gott.
Den här ölen är inte tillräckligt kall.
Den här ölen är inte kall nog.
Den här ölen har hög alkoholhalt.
Det här passet är giltigt för fem år.
Den här bussen får plats med femtio personer.
Åker den här bussen till Park Ridge?
Hur reagerade hon på nyheten?
Den här kniven är för slö för att skära med.
Den här klänningen kan se lustig ut, men jag gillar den.
Vad tycker du om den här tröjan?
Hur smakar den här soppan?
Den här datorn är bättre än den.
Adressen på det här paketet är fel.
Den här klubben har femtio medlemmar.
Jag köpte den här kameran för 35 000 yen.
Den här kameran är tillverkad i Tyskland.
Tar ni det här kortet?
Den här whiskyn är för stark.
Den här stolen är väldigt bekväm.
Var god fyll i enkäten och skicka in den till oss.
Vi har ingen snö här.
Jag hoppas att du njuter av din vistelse här.
Det här är mina skor och det här är dina.
Det är tyst här om nätterna.
Koko fortsatte att lära sig fort.
Här är din hund. Var är min?
Kan jag ställa ner den här?
För inte oväsen här.
Jag har inte sett av honom på ett tag.
Hur långt är det härifrån till Hakata?
Hur länge tar det att gå härifrån till stationen?
Vad sägs om en kopp kaffe?
Ge mig en till kopp kaffe.
Jag skulle vilja ha en till kopp kaffe.
Jag föredrar cola framför kaffe.
Hur vill du ha ditt kaffe?
Vissa gillar kaffe och andra gillar te.
Vissa tycker om kaffe och andra tycker om te.
Vissa människor gillar kaffe och andra människor gillar te.
Häng upp din kappa, tack.
Den här typen av smycken har inte mycket värde.
Ena sidan av ett mynt kallas för 'krona' och den andra kallas för 'klave'.
Ken delade rummet med sin storebror.
Vad är det Ken äter?
Ken vann över mig på schack.
Ken slog mig på schack.
Kenya blev självständigt 1963.
Tårta? Jag blev plötsligt hungrig igen.
Kate är förkyld.
Kate har tyska som huvudämne.
Kate låg ner med öppna ögon.
Vill du ha lite mer sås?
Herr Crouch, vad gör du?
Det börjar bli molnigt. Det kanske börjar regna snart.
Cuzco är en av de intressantaste platserna i världen.
Det är en vacker Kabuki docka!
Kristus tros ha utfört många underverk.
Grekiska filosofer värderade demokrati högt.
Grekerna äter också ofta fisk.
Vilket stort hus du har!
Vilket stort hus ni har!
Det regnade igår.
Han måste älska dig.
Sitt rakt.
Jag vill ha en gitarr.
Att höra är att lyda.
Ge mig nyckeln.
Torkan skadade alla skördor där.
Den stackars hunden slets bokstavligen i stycken av lejonet.
Jag blev nästan påkörd av en bil.
Var snäll och dela ut korten.
Jag tog med mig min kamera.
Det som är svårt att stå ut med är hans överdrivna artighet.
Jag har sett fram emot att få träffa dig.
Franska talas i en del av Kanada.
Det var en gång en grym konung.
Jag har coola kläder och coola solglasögon på mig.
Det tog en månad för min förkylning att gå över.
Jag ber om ursäkt för det.
Ingen orsak.
Är din mor hemma?
Tack för ditt svar.
Tack för ert svar.
Jag är utsvulten.
Far gav mig en veckas veckopeng i förskott.
Jag har blivit ombedd att informera dig om att din far har dött i en olycka.
När pappa kom hem satt jag och tittade på tv.
Vad sägs om att stanna?
Vad sägs om att sätta på en kopp te?
Du pratar så fort att jag inte förstår ett ord av vad du säger.
Jag uppskattar verkligen din vänlighet.
Kan jag få lite vatten är du snäll?
Tycker du om teatern?
Snälla låt mig få plocka upp din syster på stationen.
Diska tallrikarna är du snäll.
Låt oss hålla kontakten med varandra.
Här kommer de.
Hur mycket pengar har du?
Hur många pengar har du?
Jag är mycket glad att lära känna er.
Hur var ditt lov?
Hur var din semester?
Du då? Vill du också ha apelsinjuice?
Du då? Vill du också ha apelsinjos?
Skicka saltet.
Apelsiner innehåller mycket C-vitamin.
Vi skulle vilja beställa 18 ton olivolja.
Nederländskan är nära besläktad med tyskan.
Jag var hungrig.
Morfar pratar väldigt långsamt.
Farfar pratar väldigt långsamt.
Min farfar hör lite dåligt.
Min morfar hör lite dåligt.
Jag tar hand om min farfar.
Jag tar hand om min morfar.
Jag mår bra, tack.
Hallå där! Din baseboll hade just sönder mitt fönster.
Herregud, jag tror inte det är sant.
Låt mig se.
Jag måste ha passerat stationen medan jag tog en tupplur.
Rosorna blommar i vår gård.
Min son är längre än jag.
Eftersom han ljög straffades han.
Kaniner är besläktade med bävrar och ekorrar.
En kanin springer i trädgården.
Herr Wilson tvingade oss att upprepa meningen flera gånger.
Hur lång tid tar det att ta sig till Wien till fots?
Jag fick slut på pengar när jag var på besök i Indien.
Delfinen är ett mycket intelligent djur.
Faktum var att han till och med älskade henne.
Nu behövs inte bara ord, utan också handling.
Det är tystnad som är dyrbart nu.
Nu finns det ingen återvändo.
Jag kommer.
En hund sprang.
Hur länge har de varit här?
När kom demokrati in i existens?
Kan du säga till mig när jag ska av?
Jag vet inte precis när jag ska vara tillbaka.
Jag vet inte exakt när jag kommer att vara tillbaka.
När ska du åka till Europa?
Jag säger det hela tiden.
Kom när du vill.
Hur länge ska du vara i Japan?
Kom när ni vill.
Du kommer gilla honom så fort du fått chansen att prata med honom.
Vart fan ska du?
När fick du konsertbiljetten?
Jag träffade honom en gång.
Vi måste dra tillsammans och supa någon gång.
Hur länge har det snöat?
Italiens befolkning är hälften så stor som Japans.
En kombination av flera misstag ledde till olyckan.
En bläckfisk har tio armar.
Det är ingen bra bil, men det är en bil.
Känner du till någon bra restaurang?
Med andra ord: han är lat.
Nej, hon har aldrig blivit förälskad.
Nej, jag gick ut.
Nej, inte för mycket.
Ann spelar ofta tennis efter skolan.
Ann kommer inte till våran fest.
Va? Vad falls? Ska de inte använda sig ut av mitt förslag?
Det där är hans bil.
Det där är en pagoda.
Det är flickan som jag känner väl.
Det där är flickan som jag känner väl.
Är det en ko eller bisonoxe?
Det där är inte en gul krita.
Det där är ett bord.
Det är mitt.
Den är min.
Det där är poeten som jag träffade i Paris.
En morgon såg han en söt flicka.
Det är väldigt svårt att säga vilket land en person kommer ifrån.
En flicka ringde mig.
En tjej ringde mig.
Priset på olika maträtter varierar från vecka till vecka.
Albert, jag hoppas att du kommer stå vid mig om jag hamnar i problem.
Alice log.
I amerikansk fotboll har försvaret en specifik roll.
Amerika är ett land av invandrare.
Det finns femtio stater i Amerika.
Amerika har femtio stater.
Det liknar en anka.
Jag ska ta den jäveln.
Titta på katten.
De är för nära.
Dom säljer olika saker på den affären.
De säljer diverse varor i den affären.
Vem är den killen?
Den där röda tröjan ser bra ut på dig.
Han är bara en flyktigt bekant.
Jag lånade honom lite pengar, men han har inte betalat tillbaka dem än.
Jag lånade honom lite pengar, men har inte återbetalat dem än.
Hon kom jävligt sent.
Följ efter bilen.
Jag önskar att jag hade varit med dig då.
Den räven måste ha dödat hönan.
Håll dig undan från hunden.
Hur lång är den där bron?
Det var Herr Smith som berättade för mig hur man använde den maskinen.
Jag vill ha den väskan.
Huset är mycket gammalt. Det behöver repareras innan du säljer det.
Huset är mycket gammalt. Det behöver repareras innan ni säljer det.
Jag önskar jag kunde köpa det där huset billigt.
Ingen människa bor i byggnaden.
Ingen man bor i byggnaden.
Jag önskar att jag hade varit med henne då.
Testa den tröjan.
Du borde ha kommit med oss.
Det är en present till dig.
Du borde köpa en telefonsvarare.
Du är riktigt klusmig av dig va!
Kan du simma alls?
Du ser upptagen ut.
Är du upptagen?
Du måste hjälpa henne.
Ni måste hjälpa henne.
Känner du honom?
Pratar du japanska?
Talar du japanska?
Du har två bollar.
Du har två kulor.
Åker du med tåget eller bilen?
När brukar du vakna på morgonen?
Vem vill du prata med?
Du kan lika gärna säga det till honom i förväg.
Ni kan lika gärna säga det till honom i förväg.
Vem röstade du på i valet?
Allt du behöver göra är att vänta och se.
Du borde inte gå ut.
Du har förlorat koncentrationsförmågan.
Du påminner om en pojke som jag kände.
Känner du dem?
Känner ni dem?
Kom du med första tåget?
Du kan använda mitt skrivbord om du vill.
Har du någonsin sett en val?
Du måste gå vare sig du gillar det eller ej.
Har du någonsin varit i ett främmande land?
Ni måste hem.
Du måste hem.
Har du gjort klart din engelska läxa än?
Du får bara prata engelska.
Jag utgick ifrån att du skulle närvara på mötet.
Har du ätit färdigt frukosten än?
Du är fortfarande ung.
Allt du behöver göra är att trycka på knappen.
Vilket tåg tänker du ta?
Vet du hur man spelar schack?
Hur fick du tag på en sådan stor summa pengar?
Är du nöjd med resultatet?
Du stödjer planen, eller hur?
Du måste prata med honom angående det
Det sade du inte.
Är du för eller mot det här?
Du borde inte äta här.
Tycker du om klassisk musik?
Tror du att han är död?
Var är ditt rum?
Jag kan inte tacka nog för din vänlighet.
Om din chef "plundrar" dig betyder det att du har blivit avskedad.
Låna mig din cykel.
Vad heter du?
Vad heter du?
Jag vill ha samma ordbok som din syster.
Berätta något om ditt land.
Jag förstår inte vad du pratar om.
Jag antar att du skulle kunna ha rätt.
Jag förstår exakt hur du känner dig.
Hur skiljer sig din åsikt från hans?
Jag målade en bild åt dig.
Hur gammal är din farbror?
Hur gammal är din morbror?
Jag gav dig en bok.
Du är den sista personen jag förväntade mig att träffa här.
Du har inget att vara arg över.
Hur stor summa pengar förbrukar du?
Om du är upptagen nu kan jag ringa tillbaka till dig senare.
Du säger "dito", och det är inte detsamma som "Jag älskar dig."
Vad du har blivit lärd är fel.
Det du fick lära dig är fel.
Det ni fick lära er är fel.
Engelska kommer att ta dig en lång tid att bemästra.
Du kom in i mitt rum.
Ni kom in i mitt rum.
Ur vägen, pojk.
Jag såg mig omkring men fann ingenting.
Jag hoppas att det ska vara bra imorgon.
Jag hoppas att det är bra i morgon.
Jag älskar naturen, men jag avskyr insekter.
Vi associerar namnet Einstein med relativitetsteorin.
Tyvärr dog hon ung.
Åh, ta god tid på dig. Jag har ingen brådska.
Jag måste bege mig nu.
Aah! Min dator frös sig igen.
Vad betyder SSSR?
Vad står "PTA" för?
Två andraklassbiljetter till A är du snäll.
En 90-gradig vinkel kallas en rät vinkel.
Jag ringer dig vid sju.
Mitt plan går klockan sex.
Jag har väntat sen klockan sex och det är inte min tur än.
Ring mig klockan fyra. Jag måste ta det första tåget.
Den här målrätten är lämplig för tre.
Det började regna kraftigt för mer än tre timmar sedan.
Jag kan komma klockan tre.
Det kommer att ta tre månader för vår nya skolbyggnad att bli färdig.
Kom hit om två veckor från och med idag är du snäll.
Jag kommer tillbaka om 2 veckor.
Det går inte att säga hur långt vetenskapen kan ha nått till år 2100.
En katt dök upp från baksidan av drapperiet.
Jag måste köpa en.
Jag kommer tillbaka om en timme.
Efter klockan 11 så började gästerna att bege sig av i grupper om två och tre.
Klockan är redan elva. Det är dags att du kommer i sängs.
Kom prick klockan tio.
1,6 mil är inte en kort sträcka.
16 kilometer är inte en kort sträcka.
Kan du sänka priset till tio dollar?
Ett hundra cent blir en dollar.
Ett, tre och fem är udda tal.
"Jag är hungrig", sa den lilla vita kaninen, så de stannade och åt blomman av en stor hyasint.
"Det brinner!" skrek han.
"Är drinkarna gratis?" "Bara åt damer."
Morfar köpte den till mig.
Har du svårt med att förstå vad kvinnor och barn säger till dig?
Tror du verkligen på spöken?
Allt du behöver göra är att berätta sanningen.
Du måste inte komma hit varje dag.
Ni måste inte komma hit varje dag.
Kan du inte skilja på fantasi och verklighet?
Han är en munter kamrat.
Du är väl inte rädd för spöken?
Jag har en överraskning för dig.
Jag har en överraskning åt dig.
Jag har en överraskning åt er.
Ingen annan än du kan göra mig lycklig.
Det är upp till dig.
Du är tyst.
Var tyst.
Du ska vara tyst.
Du har förändrats.
Ni har förändrats.
Jag kan inte leva utan dig.
Jag kunde inte ta mig utanför stadion på grund av folkmassan.
Armén var tvugna att reterera.
Min bror kan komma att behöva en operation för knäskadan.
Min bror är intresserad av det man kallar popmusik.
Min bror är väldigt lång.
Direktörn kontrollerar hans män efter behag.
Jag var tvungen att överge min plan.
Polisen sa till flickorna "Är det här eran bil?"
Det var inga varningar överhuvudtaget.
Polisen hann ifatt honom.
Polisen fortsatte sin undersökning.
Polisen genomsökte det huset för att vara säkra på att de stulna skorna inte var där.
Polisen lyckades hitta brottslingen.
Jag blir hämtad.
Jag blir upphämtad.
Jag blir uppraggad.
Jag håller på att bli uppraggad.
Man trodde att valar var fiskar.
Det regnade kraftigt hela dagen.
Möt konsekvenserna.
I slutändan är det ändå talangen som räknas i musikens värld.
Han köpte den inte i alla fall.
Vi har varit gifta i fem år.
Jag sätter in tiotusen yen varje månad.
Jag sätter in tiotusen yen på banken varje månad.
Det är måndag.
Glada är de som känner till värdet av hälsa.
Hunden bet mig i handen.
En hund skäller.
Har du matat hunden än?
Hunden har bitit hål på min ärm.
Kan du finna den?
Kan du hitta den?
Så långt ögat kunde se var marken täckt med snö.
En vis man drar nytta ut av sina mistag.
Jag letar efter min nyckel.
Lycka till.
Ryck upp dig!
Ryck upp er!
Var bor du nu?
Var bor ni nu?
Verklighet och fantasi är svåra att skilja på.
Det här är året av information, och datorer spelar en ökande viktig roll i vårt vardagliga liv.
Lättare sagt än gjort.
Jag undrar om det finns någon mening i att lägga in ordspråk i engelskan?
Andas han?
Döm inte andra efter dig själv.
Lås dörren!
Sjön hade frusit till, så vi gick över isen.
Det kommer att regna den här eftermiddagen.
Efter oss syndafloden.
Var snäll och stäng dörren efter dig.
Missförstå mig ej, vi gör inga löften.
Du skall observera trafikreglerna.
Anledningen till trafikolyckan rapporterades av polisen.
Jag hittade en bebis fågel när jag gick i parken.
Öppna din mun.
Öppna munnen.
Du pratar för mycket.
Kvinnan som sitter där borta är hans nuvarande fru.
Vem är flickan som står där borta?
Gör vad du vill.
Du får prata hur mycket du vill.
Vilket märke gillar du?
Nyfikenhet dödade katten.
Som tur är blev ingen blöt.
Som tur är var vädret bra.
Lyckan log mot honom.
Ett mynt ramlade ut ur hans ficka.
En kopp te, tack.
Vad sägs om en kopp te?
Fundera på det.
De som inte önskar gå behöver inte det.
Jag ger upp.
Kasta inte in handduken.
Några är dyra medan andra är väldigt billiga.
Förenta nationerna är en internationell organisation.
Jag är upptagen nu.
Tiden är mogen för en drastisk förändring.
Nu eller aldrig.
Får jag titta på tv nu?
Jag är inte mannen som du en gång kännde mig som.
Jag känner inte för att äta just nu.
Om jag var rik så skulle jag åka utomlands.
Om jag vore rik, skulle jag åka utomlands.
Vad är populärt nu?
Vad är inne nu?
Vad är på modet nu?
Vad är klockan? Min klocka går fel.
Jag kan inte komma av arbetet nu.
Till slutet av veckan.
När gick du upp imorse?
Kom ihåg att följa med mig och fiska på söndag.
Jag tror inte att det kommer att regna i eftermiddag.
Är du ledig i eftermiddag?
Du måste intressera dig för aktuella händelser.
Du kommer inte att finna så många nyheter i dagens nyhetstidning.
I morse klarnade det.
Låt oss stoppa här.
Vi stannar här.
Jag är inte säker på att vi kommer kunna få tag på biljetter ikväll.
Det är galet varmt idag.
Vill du inte simma idag?
Vill ni inte simma idag?
Jag känner inte för att äta någonting idag.
Det ska bli kallare och snöa senare idag.
Jag har inga lektioner idag.
Jag har matteläxa idag.
Jag vill inte träffa någon i dag.
Skrev du något i din dagbok idag?
Jag är ganska trött idag.
Det här är den kallaste vintern som vi har haft på trettio år.
Vad sägs om att spela schack i kväll?
Vi väntar främmande i kväll.
Jag ringer honom ikväll.
Vad ska du göra ikväll?
Månen är mycket vacker i kväll.
Han är i tjänst inatt.
Problemet med honom är att han är lat.
Problemet är att vi inte har någonstans att vara ikväll.
Vi har inget socker.
Håll bollen i rullning.
De som styr mest gör minst ljud ifrån sig.
En färsk undersökning visar att antalet rökare minskar.
Jag minns den första gången.
Först visste jag inte vad jag skulle göra.
Först visste jag inte vad jag skulle ta mig till.
Först trodde jag att han var lärare, men det var han inte.
En man vars fru är död kallas för en änkling.
Den finansiella situationen förvärras vecka för vecka.
Hela dagen var min pappa på dåligt humör för att han tappat bort sin plånbok.
Lägg inte plånboken på elementet.
Lägg inte plånboken ovanpå elementet.
Har du skrivit klart din uppsats?
Jag har inte ätit något sedan i går.
Det var söndag i går, inte lördag.
I går var det söndag, inte lördag.
Igår var han väldigt sjuk men idag mår han mycket bättre.
Det var hans bil, inte min, som gick sönder igår.
Stålproduktion nådde uppskattat 100 miljoner ton förra året.
Jag är trött eftersom jag var tvungen att plugga inför ett prov igår natt.
Vad gjorde du i går kväll?
Tjuvar bröt sig in i mitt hus i går kväll.
Tallriken slank från hennes hand och krashade ner i golvet.
Jag brukar diska.
Jag måste ta ett paraply med mig.
Repet gick av medan vi besteg berget.
Skulle du vilja följa med på en promenad?
Jag fruktar det.
Jag står inte ut att bli störd i mitt arbete.
Arbetsnarkomaner ser semesterdagar som slöseri med tid.
Arbetsnarkomaner ser semester som tidsslöseri.
Du gillar visst inte sashimi?
Jag är på väg till min systers bröllop.
Sluta bete dig som ett barn.
Två läsk till barnen och en kaffe, tack.
Stick härifrån, ungjävlar!
Det finns en park i centrum.
Hans utställning på stadsmuséet tilltalade mig inte alls.
Förutom borgmästaren var många andra förnäma gäster närvarande.
Tankar uttrycks genom ord.
Tankar uttrycks med hjälp av ord.
Hisaos ansikte var likblekt.
Jag lagade kvällsmat.
Tio år har gått sedan jag kom hit.
Det har gått tio år sedan jag kom hit.
Det tog mig tre dagar att läsa den här boken.
Jag fick reda på det av en ren händelse.
Måste jag hålla ett tal?
Jag försörjer min familj.
Ser du efter barnen medan jag är ute?
Ken läste när jag kom hem.
Det här skrivbordet som jag köpte igår är väldigt stort.
Jag tar det.
Om hon bara hade vetat att jag var i Tokyo, skulle hon ha hälsat på mig.
Det är allt jag känner till om honom.
När jag besökte deras lägenhet var paret precis i ett gräl.
Jag erkänner att jag är slarvig.
Det var min tur att städa rummet.
Mannen som jag besökte var Mr Doi.
Vänta här tills jag kommer tillbaka.
Han sa ingenting medan jag talade.
Det fanns ingen kvar utom mig.
Vi iakttog honom tills han var utom synhåll.
Varför följer du inte med oss till festen?
Vårt lag besegrade motståndaren med 5-4.
Vår engelsklärare lägger vikt vid uttalet.
Vår skola är femton år gammal.
Vårt lov kommer snart att nå sitt slut.
Vår plan kommer att fungera bra.
Vår bil är tre år äldre än er.
Vår bil är tre år äldre än din.
Vår bil är tre år äldre än era.
Vår bil är tre år äldre än dina.
Jag kan inte komma på något annat sätt att få honom att acceptera vårt förslag.
Vi försöker.
Vi är människor.
Vi är hans söner.
Fast att vi väntade till tio dök Bill aldrig upp.
Vi vann matchen med 10 mot 4
Vi är tacksamma för er vänlighet.
Vi är tacksamma för din vänlighet.
Vi körde för snabbt för att njuta ut av det vacka landskapet.
Vi har för många lektioner.
Vi är inte amerikaner.
Vi kommer alltid att vara tillsammans.
Vi talar i Australiens ungdomars vägnar.
Vi hade roligt på stranden igår.
Vi genomförde vår utredning med största noggrannhet.
Vi måste ta itu med det här problemet.
Vi fick aldrig någon tydlig förklaring på mysteriet.
Vi såg barnet kliva på bussen.
Vi såg barnet stiga på bussen.
Vi satt mitt i rummet.
Vi trodde att det var ett flygande tefat.
Vi visste inte vad vi skulle göra.
Vi hade väldigt kul.
Vi måste försvara vårt land till varje pris.
Vi använder ätpinnar istället för kniv och gaffel.
Vi lärde oss ryska istället för franska.
Vi flög från London till New York.
Vi såg något vitt i mörkret.
Vi bor nära stationen.
Vi är alla överens med er.
Vi är alla överens med dig.
Vi flyttade våra väskor för att ge plats för den gamla damen att sitta ner.
Vi gick på picnic till kullen.
Vi är rädda.
Vi lär oss om antikens Rom och Grekland.
Vi njöt av att simma i sjön.
Vi lekte ofta mamma pappa barn i parken.
Vi tillbringade en natt i en fjällstuga.
Vi åker och fiskar då och då.
Vi lyssnar med öronen.
Vi satte oss i bilen.
Vi prövar en helt ny metod.
Vi är mer eller mindre själviska.
Vi föddes på samma dag.
Vi var fattiga, men glada.
Vi sover vanligtvis i det här rummet.
Vi spelade baseball.
Jag satte upp en liten koja i trädgården.
Vi dekorerade rummet själva.
Jag är typen som skyr risker som pesten.
Jag har varit bekant med henne i över 20 år.
Jag har känt henne i över 20 år.
Den här boken är för mig vad Bibeln är för dig.
Det är svårt för mig.
Jag har en vän vars far är kapten på ett stort skepp.
Jag gillar inte modern jazz.
Jag har två utländska vänner.
Jag antar att du beredd på att ta risken.
Jag antar att du är beredd att ta risken.
För min del föredrar jag öl framför whisky.
Jag bjuder.
Min klass består av fyrtio studenter.
Kommer du ihåg mig?
Mitt skägg växer snabbt.
Min åsikt skiljer sig från din.
Min engelska är allt men inte bra.
Min engelska är allt utom bra.
Mitt sommarlov är över.
Mitt hus ligger tio minuters gångväg från stationen.
Mina skor måste lagas.
Han är min bror.
Min bror bor i en liten by.
Min bror är bra på tennis.
Min storebror är lärare.
Min bror bor i Tokyo.
Min bror anländer imorgon bitti.
Min hund låtsas ofta sova.
Min hund är vit.
Kan du höra mig?
Kan ni höra mig?
Min lycka beror på dig.
Min åsikt skiljer sig från din.
Båda mina systrar är gifta.
Min cykel behöver lagas.
Mitt uppslagsverk är väldigt användbart.
Min ordbok är mycket användbar.
Det är något fel på min bil.
Min bil håller på att bli reparerad nu.
Min bil är stor nog för fem personer.
Jag hittar inte min portfölj.
Mitt huvudämne är europeisk medeltidshistoria.
Så vitt jag vet håller de alltid sina löften.
Min bror har aldrig bestigit Mt Fuji.
Min bror är lika lång som jag.
Min bror kan springa lika fort som jag kan.
Min bror måste skriva en tentamen.
Mitt hår är längst i klassen.
Min far varken röker eller dricker.
Min far är duktig på att simma.
Mitt rum är mycket litet.
Mitt rum vetter mot öst.
Min mor tar en tupplur varje eftermiddag.
Jag är längre.
Min dröm är fortfarande bara en dröm.
Min väckarklocka ringde inte i morse.
Jag äter upp min hatt om min kandidat inte vinner valet.
Jag hoppas att din förkylning går över snart.
Jag gillar österrikisk musik.
Jag tycker om österrikisk musik.
Jag börjar så sakta tycka om Ken.
Jag spelade fotboll igår.
Jag är ansvarig för hans beteende.
Jag beställde nya möbler.
Jag lärde mig att cykla när jag var sex år gammal.
Jag gav dem ett tusen yen var.
Jag tar ett bad varannan dag.
Jag har läst engelska i fyra år.
Jag har studerat engelska i fyra år.
Jag har varit här sedan klockan fem.
Jag stannar här till i övermorgon.
Jag håller inte med dig.
Jag tackar dig.
Jag tackar er.
Jag skulle vilja att du betalar i förskott.
Jag är dubbelt så gammal som du.
Jag tänker på dig hela tiden.
Jag kommer aldrig att glömma din vänlighet.
Jag kan inte besvara din fråga.
Jag uppskattar vår vänskap mycket.
Jag tycker att den sociala sidan är intressant i den nyhetstidningen.
Jag skaffade en ny högtalare i den affären.
Jag bor i en lägenhet.
Jag bor i lägenhet.
Jag åkte till Europa via USA.
Jag gick och lade mig lite senare än vanligt.
Jag har alltid en ordbok nära till hands.
Jag blev bortförd av utomjordingar.
Jag blev bortförd av rymdvarelser.
Jag blev kidnappad av rymdvarelser.
Jag blev kidnappad av utomjordingar.
Jag har aldrig varit hemma hos min farbror.
Jag har aldrig varit hemma hos min morbror.
Jag har precis varit på stationen för att vinka av min farbror.
Jag har precis varit på stationen för att vinka av min morbror.
Jag tycker bättre om roliga filmer.
Jag bor intill leksaksaffären.
Jag är inte så förtjust i grönt te.
Jag gillar te.
Jag tycker om te.
Min mor brukade läsa sagor för mig.
Jag tenderar till att dra till mig förkylningar.
Jag kan spela gitarr.
Jag studerade en stund i morse.
Jag pluggade en stund i morse.
Jag gillar inte klassisk musik.
Jag har bott här
Jag letar efter en man som ska bo här.
Jag har hållit på att skriva det här manuskriptet i ett år.
Jag är nöjd med de här skorna.
Jag vet inte vad det här ordet betyder.
Jag tror inte på att det finns någon ond person i denna värld.
Jag skulle vilja simma i den här floden.
Jag böjer mig inte en millimeter i den här frågan.
Det tog mig en halvtimme att lösa det här problemet.
Jag har ingen aning om hur man spelar golf.
Jag yrkar att vi godkänner förslaget och att åtgärder vidtas så fort som möjligt.
Jag skakade hand med Jane.
Jag är inte det minsta förvånad.
För länge sedan besökte jag Kanada.
Jag har varit upptagen.
Jag blev blöt ända in på skinnet.
Jag tror det.
Jag hade ingenting att göra med gruppen.
Jag gillar varken den ena eller den andra kakan.
Det visste jag inte.
Jag visade dem hur man gör det.
Jag visade för dem hur man gör.
Jag funderade på planen.
Jag kom enbart för att ge besked om faktumet.
Jag såg bilen köra på en man.
Jag står inte ut med oljudet längre.
Jag minns mannens ansikte men jag kommer ej ihåg hans namn.
Jag har inget med brottet att göra.
Jag sträckte ut handen mot boken.
Jag har inte läst boken och inte vill jag göra det heller.
Jag gick upp tidigt för att hinna med tåget.
Jag kan sjunga det på engelska.
Jag använder det.
Jag kan inte göra något sånt.
Jag har massor av kameror.
Jag har bara en önskan.
Jag stod och väntade på en buss.
Jag kan inte röka.
Jag pluggade i kanske två timmar.
Jag börjar komma ihåg det.
Jag vann över honom på schack.
Jag slog honom på schack.
Jag har en bok om fiske.
Jag är dålig på tennis.
Jag tycker om tennis.
Jag känner tjejen som spelar tennis.
Han spelade tennis.
Jag klarar av att försörja min familj.
Ibland känner jag mig ledsen.
Var är jag?
Jag gillar båda.
Jag hade en väldigt hög feber.
Jag gillade Tony.
Jag vet inte hur man köper en biljett.
Jag vill ha en Toyota.
Jag skulle vilja bo i New York.
Jag har en katt och en hund. Katten är svart och hunden är vit.
Jag såg henne på festen.
Jag har varit i Paris.
Jag kan inte läsa franska, inte heller kan jag tala det.
Jag kan inte läsa franska, och ännu mindre tala det.
Jag har en penna.
Jag avbröt min hotelreservation.
Jag har redan gjort det.
Jag har redan gjort det.
Jag behöver inte gå till doktorn längre. Jag mår mycket bättre.
Jag måste bege mig nu.
Jag kommer inte att träffa henne igen.
Jag gillar att ha mycket att göra.
Jag brukade åka skidor på vintrarna.
Jag blir ofta förkyld.
Jag älskar rock.
Jag åkte ända till London med bil.
Jag har klättrat upp för berget Aso.
Jag är en doktor.
Jag köpte en bok.
Jag går till biblioteket två till tre gånger om veckan.
Jag går till biblioteket två eller tre gånger i veckan.
Jag går till biblioteket två till tre gånger per vecka.
Jag är van vid att jobba hårt.
Jag är van vid att arbeta hårt.
Jag har bestämt mig för att gå i pension.
Jag hade tur.
Jag ska sluta röka för gott.
Jag kan simma.
Jag gillar engelska, men jag är inte så bra på att tala det.
Jag vill inte sjunga, för jag är tondöv.
Jag vet inte vad klockan är.
Jag har mitt eget sovrum hemma.
Jag sköt upp hushållsarbetet några timmar.
Jag sköt upp mitt hushållsarbete några timmar.
Jag sköt på mitt hushållsarbete några timmar.
Jag har många blommor. Några är röda och andra är gula.
Jag gillar att ta mitt block och min penna och åka till kusten för att skissa.
Jag presenterade mig på mötet.
Jag ångrar att jag var så lat under min skoltid.
Jag kan knappt se utan mina glasögon.
Det kändes som om mitt ansikte brann.
Får jag gå hem?
Jag åt snabbt upp min lunch.
Jag vill dricka mjölk.
Jag hade en intressant konversation med min granne.
Jag vill be dig om en tjänst.
Jag vill att du läser det här engelska brevet.
Jag känner din bror väl.
Jag kanske skriver ett brev åt dig.
Jag spelade tennis med min bror.
Jag är ekonomiskt självständig från mina föräldrar.
Jag åker till Hiroshima tre gånger i månaden.
Jag kännde igen henne stunden jag såg henne.
Jag såg en gammal vän.
Jag gillar att gå en tur i parken.
Jag har inget emot det.
Jag vill dricka en kopp te.
Jag råder dig att inte åka.
Jag gick inte, utan stannade hemma.
Jag är upptagen med maten för tillfället.
Aldrig hade jag sett en sådan fridfull syn.
Jag har läst några hundratals böcker.
Nu är jag på flygplatsen.
Jag kommer inte på hans namn just nu.
Jag brukar inte dricka kaffe utan socker.
Jag såg honom igen.
Jag tror att ärligheten kommer att vinna i slutändan.
Det var inte förrän igår jag fick nyheterna.
Jag lämnade in ett papper igår.
Jag steg upp tidigt igår.
Jag läste ut boken i går kväll.
Jag luktar med näsan.
Jag är älskad av mina föräldrar.
Jag tänker skriva om våra parker och berg.
Jag har varit hos tandläkaren.
Jag vill ha ett eget rum.
Jag höll i festen på egen bekostnad.
Jag vill tro att jag vet vad jag pratar om.
Jag kan bara tala för mig själv.
Jag gjorde det mot min vilja.
Jag minns huset som jag växte upp i.
Jag trodde inte mina ögon.
Jag gick hemifrån vid sju.
Jag ska köpa en bil.
Jag har tillräckligt med pengar för att köpa en bil.
Jag gav tillbaka kniven som jag hade lånat.
Jag har inte tid att göra mina läxor.
Jag har aldrig blivit kär i någon tjej.
I framtiden vill jag bli en TV-presentatör.
Jag har lite pengar.
Jag är inte ett dugg trött.
Jag fick syn på pojken.
Jag var född och uppfostrad i Matsuyama.
Jag kan simma bra.
Jag diskar.
Jag försov mig.
Jag har byggt ett nytt hus.
Jag byggde ett nytt hus.
Jag såg på när den röda solen gick ner i väst.
Jag förlorade henne ur sikte i folksamlingen.
Jag gillar att läsa deckaren.
Jag gillar att simma.
Jag tycker om att simma.
Jag tycker om simning.
Jag tycker om att simma, men inte här.
Jag ämnade att lyckas, men kunde inte.
Jag avskyr politik.
Jag har inte sett henne sen förra månaden.
Jag är lärare.
Jag fick min son till att träffa doktorn.
Jag är hälsosam.
Mitt huvudämne på universitetet var kemi.
Jag representerade mitt universitet på konferansen.
Jag gick längs huvudgatan.
Jag är hungrig för jag har inte ätit lunch.
Jag träffade Fred på gatan.
Jag kommer att åka oavsett väder.
Jag väntar på att affärens ska öppna.
Jag gillar vinter.
Jag tog hans närvaro för givet.
Jag stannar här tillsvidare.
Han kan varken läsa eller skriva.
Jag bor i Japan.
Jag återvände till Japan.
Jag är japan, men du är amerikan.
Jag är gravid.
Jag har ingen katt.
Jag släppte in katten i mitt rum.
Jag arbetade på en bondgård.
Jag har en svår smärta i ryggen.
Jag såg en vit hund hoppa över staketet.
Jag misstänkte att han ljög, men det kom inte som en överraskning.
Jag är förvånad att han antog erbjudandet.
Jag är förvånad att han accepterade erbjudandet.
Jag vet inte vad han har råkat ut för.
Jag vet inte vad som har hänt med honom.
Jag vet var han bor. Men det är en hemlighet.
Jag är skyldig honom 100 yen.
Jag trodde att han var en doktor.
Jag frågade vem han var.
Jag rådde honom att komma tillbaka omedelbart.
Jag hittade en fin lägenhet åt honom.
Jag varnade honom för faran.
Jag hittade ett jobb åt honom.
Jag förklarade det för honom, bara för att förvirra honom.
Jag frågade honom vad han hette.
Jag vill veta orsaken till hans frånvaro.
Jag kunde inte förstå något ut av vad han sa.
Jag observerade att hans händer var ostadiga.
Jag fick ett brev som informerade mig om hans ankomst.
Jag fick ett brev som underrättade mig om hans ankomst.
Jag drömde om honom.
Jag är hans vän och kommer så förbli.
Jag åkte till flygplatsen för att träffa honom.
Jag åkte till flygplatsen för att möta upp honom.
Jag fick veta att det var svårt för henne att lösa det problemet.
Jag såg henne simma.
Jag hjälpte henne med att hänga upp bilden på väggen.
Jag vet att hon har varit upptagen.
Ju mer jag lyssnar på henne, desto mindre gillar jag henne.
Jag vill komma i kontakt med henne.
Jag sa till henne att kvickt göra klart rapporten.
Jag ämnade ringa henne, men jag glömde att göra det.
Jag försökte ge henne en gåta.
Jag älskar henne.
Jag var oförmögen att titta henne i ansiktet.
Jag är orolig för hennes hälsa.
Jag gissade att hon var fyrtio.
Jag tror på hennes berättelse.
Jag föreslog honom att hon skulle bli inbjuden till festen.
Jag tittade på henne.
Jag kunde hjälpa henne.
Jag föredrar komedier framför tragedier.
Jag var trött.
Även om jag var trött så försökte jag mitt bästa.
Jag var väldigt trött, så jag gick och la mig tidigt.
Jag åkte flygplan till Kyushu.
Jag åkte till Kyushu med flygplan.
Jag vill lära mig standardengelska.
Jag gick inte på grund av sjukdom.
Jag tror att jag har råkat på en förkylning.
Jag ringde inte honom eftersom jag hade en förkylning.
Jag sprang till min mamma.
Jag ska spela fotboll efter skolan.
Jag är upptagen.
Jag sålde en bok.
Jag är riktigt oroad över din framtid.
Jag använder det varenda dag.
Jag promenerar i skogen varje dag.
Jag springer varje dag.
Jag joggar varje dag.
Jag är rädd för vilda djur.
Jag kände mig smått illamående.
Jag var kolugn.
Jag vill studera utomlands.
Jag vill plugga utomlands.
Jag sprang så snabbt jag kunde för att hinna med tåget.
Jag gick också.
Jag önskar att jag kunde simma lika långt som han.
Tar du mig för fyrtio? Du missar rejält!
Titta på mig.
Jag har många vänner som hjälper mig.
Jag önskar att jag hade ett eget rum.
Jag önskar att jag hade ett rum för mig själv.
När vi kom hem hade solen gått ner helt och hållet.
Var snäll och ge oss två knivar och fyra gafflar.
Vår fotbollsmatch kommer att skjutas upp.
Vår lärare skrattar sällan.
Vi ska mötas vid sju.
Vi hyrde en lägenhet.
Vi tillbringade en utmärkt semester i Sverige.
Vi förknippar namnet Darwin med evolutionsteorin.
Vi råkade befinna oss på samma buss.
Vi lyckades simma över ån.
Vi såg inget konstigt.
Vi träffas här en gång i månaden.
Vi såg många skepp i hamnen.
Vi kan inte vara utan vatten ens för en dag.
Vi klev upp tidigt så att vi kunde se soluppgången.
Vi steg upp tidigt så att vi kunde se soluppgången.
Vi tipsade dom om att börja tidigt.
Vi hoppas på fred.
Rita ett streck på ditt papper.
Jag försökte skriva med min vänstra hand.
Jag är rädd att jag inte kommer att vara ledig förrän examinationen är slut.
Det blev oavgjort.
Matchen kan ha skjutits upp till nästa vecka.
Vi blir tvungna att skjuta upp matchen till nästa söndag.
Jag har en fruktansvärd tandvärk.
Har du borstat tänderna?
Jag måste träffa en tandläkare.
Jag kan inte komma på någon bra ursäkt till varför jag är sen till tandläkaren.
Tandläkaren drog ut hennes dåliga tand.
Orsaken till olyckan är okänd.
Han reflekterade över hur snabbt tiden går.
Tiden flyger.
Tiden rusar.
Han sprang för att komma i tid.
En dator är inte mer levande än vad en klocka är.
Jag tappade bort klockan.
Säg vad vi ska göra härnäst.
Till jul har vi känt varandra i tre år
Hur långt ifrån ligger nästa bensinstation?
Jag blev tvungen att vänta i tjugo minuter på nästa bus.
Jag ska av nästa station.
Jag ser fram emot att få träffa dig nästa söndag.
Var skulle du vilja åka nästa söndag?
Hur dags går nästa tåg till Tokyo?
Han gräver sin egen grav.
Det läker av sig själv.
Ställ undan cykeln.
Jag känner mig som en annan person.
Jag vill hålla mitt rum så prydligt som möjligt.
Låt mig betala min del.
Jag trodde knappt mina ögon.
Gör gott mot dem som hatar er.
Gören gott mot dem som hata eder.
Ingenting saknas.
Jag håller inte med.
Jag tog mig friheten att ringa henne.
Ditt svar på frågan visade sig vara fel.
Faktum är att han inte håller med mig.
Faktum är att hon läste inte ens brevet.
Ärligt talat har jag redan sett den filmen.
Sanningen att säga, led änkan av magcancer.
Om jag ska säga sanningen minns jag ingenting jag sa i går.
Experimentet var lyckat.
Faktum är att han är troende.
Det hände egentligen inte.
Jag önskar att jag hade en bil.
Titta på pojken bredvid bilen.
Kör försiktigt.
Jag glömde mina bilnycklar.
Vad har du gjort angående reperationen av bilen?
Bilen körde in i ett skyddsräcke.
Få jag låna din bil?
Troligt är att inget språk fullständigt saknar lånord.
Ung som han är kan han arbeta hela dagen lång.
Du är bara ung en gång.
En ung flicka satt vid ratten.
Vem spelar huvudrollen?
Jag ringer min man.
Jag har inte så mycket pengar med mig.
Det är nödvändigt att bekämpa AIDS med vilket vapen vi nu än behöver!
Släpp inte taget.
Brevets innehåll var hemligt.
Påminn att posta breven är du snäll.
Får jag hjälpa?
På grund av den dåliga skörden har vetepriset gått upp de senaste sex månaderna.
Religion är ett opium för folket.
Löven ändrar färg i höst.
Det var snällt av dig att hjälpa mig med läxan.
Det är dags att åka.
Det är dags att gå.
Släpp ut mig!
Var är utgången?
Skadorna från översvämningen räknas bli tio miljoner dollar.
Föräldrarna var förtjusta av hennes skönhet.
Jag ska göra mitt bästa.
Vänta på din tur.
Det är svårt för en nybörjare att uppskatta vindsurfing.
Det var varmt, och fuktigt till yttermera visso.
Det var varmt och dessutom fuktigt.
Det är för varmt.
Snälla hjälp mig.
Hon ville veta om fotografen kunde ta bort hatten från bilden.
Var har bildats i såret.
Pilla inte på såret.
Låt inte din fantasi springa iväg.
Vi är säkra på vår vinst.
Jag förväntar mig en tunnelbanestation här i framtiden.
Det är omöjligt att veta vad som kommer att hända i framtiden.
Den är för liten.
Det är för litet.
Det lilla födelsemärket tog ingenting ifrån hennes skönhet
Sluta reta mig.
Tjejer kom in, den ena efter den andra.
Flickor kom in, den ena efter den andra.
Flickan var snäll och berättade vägen till museet.
Flickan var alldelles utom av sig av sorg.
En pojke sprang iväg med lite pengar.
De lade ut mattan på golvet.
Tack så mycket för att ni bjöd in mig.
Tack så mycket för att du bjöd in mig.
Får jag låna ditt suddgummi?
Var är rulltrappan upp?
Senatorn anklagade mig för att ha förvrängt datan.
Vill du ha lift?
Vill du ha skjuts?
Det är inget skämt.
Du måste skämta!
Du bör alltid tänka innan du talar.
Man bör alltid tänka innan man talar.
Han hade i arbetet kommit i kontakt med några utlänningar.
Ät så mycket du vill.
Du får inte läsa, medan du äter.
Om man äter för mycket blir man tjock.
Om du äter för mycket kommer du att bli tjock.
Efter måltiden frågade jag efter räkningen.
Det är viktigt att följa en sträng diet.
Det är otroligt.
Signalen blev grön.
Trafikljuset slog om till rött.
Jag har nariga läppar.
Det tog hela kvällen.
Domaren utgav honom som vinnare.
Oro gjorde mig sömnlös igår natt.
Jag ska köpa en ny.
Hur är den nya ledaren?
Jag behöver en ny cykel.
Släpp in lite frisk luft.
Var är tidningen?
Enligt tidningen ska det snöa imorgon.
Det stod i tidningen att ännu ett krig har brutit ut i Afrika.
Allt var fortfarande i skogen.
Jag är ledsen, vi har inga vaccin.
Tyvärr, jag har ingen aning.
Det är svårt att skilja sanning från lögn.
Du dödar mig långsamt.
Mari och Maki är systrar.
I begynnelsen skapade Gud himmel och jord.
Gud skapade världen på sex dagar.
Föräldrar älskar sina barn.
Jag bröt av min tumnagel.
Det är iskallt.
Har du någon legitimation?
Man lär sig ut av erfarenheter.
Ju mer vi har desto mer vill vi ha.
Det är nödvändigt för oss att sova gott.
Skämtar du?
Peka inte på andra.
Det är oartigt att peka på folk.
Folk älskar frihet.
Människorna skrattade tills hon sa "Brinn!".
Förr trodde man att bara människor kunde använda språk.
Var rädd om dina möten med andra för du vet aldrig om du bara möter personen en gång om livet.
Om inte människan tar hand om miljön kanske miljön eliminerar mänskligheten.
Utan vatten så skulle vi snart dö.
Det är omöjligt att leva utan vatten.
Vatten, tack.
Lägg till vatten och blanda ihop det till en mjuk deg.
Du borde verkligen inte dricka kranvattnet.
Du måste få tillräckligt med sömn.
Det finns mer än 4000 språk i världen.
Ingen kan förneka faktumet att världsekonomin kretsar kring den amerikanska ekonomin.
Vi måste avsluta det här arbetet till varje pris.
Vare sig du lyckas eller inte beror på dina egna ansträngningar.
Om någon är politiker är det han.
Det är mycket ovanligare för en person att vara politiskt medveten än att vara politiskt aktiv.
Stjärnorna blinkade på himlen.
Ibland är det svårt att skilja rätt från fel.
Gör det som du tycker är rätt.
En nyfödd baby är benägen att bli sjuk.
Produktionen har börjat avta.
Många av eleverna var trötta.
Studenterna delade in sig i tre grupper.
Lärarens elever ser upp till honom.
Det finns inget annat att göra än att vänta på att platserna blir lediga.
Jag skulle vilja byta plats.
Det var en gång en stor konung som bodde i Grekland.
Det var en gång en fattig man och en rik kvinna.
Tvål har förmågan att få bort smuts.
Kolet glöd i elden.
Har du namngett din nyfödda bäbis?
Ett spädbarn sover i vaggan.
Spädbarnet log mot mig.
Barnet slutade gråta.
En bebis är inkapabel ut av att ta hand om sig själv.
Underskottet har minskat lite i taget.
Du kan köpa frimärken på vilket postkontor som helst.
Ni kan köpa frimärken på vilket postkontor som helst.
Man kan köpa frimärken på vilket postkontor som helst.
Biljetterna är slutsålda.
På grund av snön så missade jag tåget.
Matchen blev fördröjd på grund ut av snö.
Det fortsatte att snöa i fyra dagar.
Jag är helt säker!
Senaste gången var det en naturlig födelse.
Varorna som beställdes från England förra månaden har inte anlänt än.
Vad gjorde du förra söndagen?
Fram tills förra veckan hade jag inte fått något svar.
Här kommer vår lärare.
Läraren tolkade meningen åt oss.
De fortsatte att prata, till och med efter att läraren kom in.
Där kommer vår lärare.
Varför frågar du inte din lärare om råd?
Läraren underströk vikten av att föra anteckningar.
Läraren öppnade lådan och tog ut en boll.
Jag gjorde ett försök att simma över floden.
Jag vill ha fläkten.
Skeppet sjunker.
Valets resultat kommer snart att bli analyserad.
Valresultatet kommer snart att analyseras.
Du stötte på honom tidigare, eller hur?
Ni stötte på honom tidigare, eller hur?
Den förra hyresgästen skötte lägenheten utmärkt.
Visst är det vackert väder?
All kunskap är inte till godo.
Vi är femton, allt som allt.
Hela nationen sörjde hjältens död.
Mormor bar bordet själv.
Farmor bar bordet själv.
Kom hem tidigt, Bill.
Titta inte ut genom fönstret.
Öppna fönstret.
Stäng fönstret.
Skulle du kunna slå in den som en gåva?
Hennes söner har åkt till Tokyo.
Sonen ställde en fråga till hans mor.
Se upp var du går.
Spring fort, annars kommer du för sent till skolan!
Lätt gånget lätt förgånget.
Inte en människa syntes till i byn.
Det finns en sjö öster om byn.
Jag kan inte tänka mig något annat.
Han har bara en tröja för resten av dom är på tvätt.
De andra barnen skrattade.
Man ska inte göra sig lustig över andra.
Många utlänningar pratar bra japanska.
Många unga i Japan äter bröd till frukost.
Tillåt inte dig själv att bli tjock.
Stilla Havet är det största havet i världen.
Solen gör jorden varm och ljus.
Solen går upp i öst och ner i väst.
Har du gått ner i vikt?
Jag kan inte direkt säga att jag är glad över min pensionering.
Där är en katt i köket.
Det är en katt i köket.
Det finns en katt i köket.
Vad du har växt!
Det är för högt.
Ett stort djur sprang iväg från zooet.
Det tunga regnet förhindrade mig från att komma ut.
Luftföroreningar är ett allvarligt globalt problem.
Massorna reste sig mot diktatorn.
Vi har large, medium och small. Vilken storlek vill du ha?
Vi har large, medium och small. Vilken storlek vill ni ha?
Att bo i en storstad har många fördelar.
Presidenten är för närvarande i Miami.
Sedan jag återhämtade mig från min allvarliga sjukdom ter sig hela skapelsen vacker för mig.
När bröt andra världskriget ut?
Vem springer snabbast i din klass?
Vem upptäckte Amerika?
Någon har stulit alla mina pengar.
Jag hörde någon skrika.
Jag behöver någon.
Vem kan utföra det här arbetet?
Vem skrev det här brevet?
Vet du vem som har skrivit den här romanen?
Finns det någon som kan uttala det här ordet?
Vem tycker inte så?
Är någon hemma?
Kan någon annan svara?
Vem vet?
Det finns inget ont som inte har något gott med sig.
Hur firade du din födelsedag?
Männen gick för att jaga lejon.
Pojkar härmar ofta sina idrottshjältar.
Både pojkar och flickor borde studera hemkunskap.
Vem vet inte?
Kunskap är makt.
Jorden är ingen stjärna, utan en planet.
Inget är så hemskt som en jordbävning.
Dammen har torkat ut.
Det var just likt honom att komma för sent.
Du är sen.
Du är inte i tid.
Vem är den där kvinnan i brun jacka?
Släpp in mig.
Kan du räkna till tio på kinesiska?
Försiktig som han var gjorde han ett oväntat misstag.
Lyssna noga är du snäll.
Jag är ingen morgonmänniska.
Frukosten är färdig.
Frukost är en smörgåsbord.
Har du någonsin varit på Koreahalvön?
Gå upp tidigt på morgonen.
Det är skönt att stiga upp tidigt.
Vi tappade bort tornet när vi gick in i byn.
Publiken bestod mest ut av elever.
Publiken såg uttråkad ut.
Jag väntade inte länge förän han dök upp.
Den långa resan förvärrade hennes skada.
Fåglar sjunger.
Fåglar flyger.
Fåglarna lägger ägg.
Det är ovanligt.
Vilken lägenhet som helst duger så länge hyran är rimlig.
Det ligger affärer längs gatan.
Varför inte ansöka om jobbet som tolk?
Lägg inte dina grejer i gången.
Där är vackra blommor här och där i trädgården.
Med små steg började rosbuskens knoppar blomma.
Kan du säga namnet på alla träd i trädgården?
Trädgårdsmästaren planterade en ros mitt i trädgården.
Min bror måste ha skrivit det här brevet.
Min bror vågade ej att simma över floden.
Ge inte upp!
Lera är en grundläggande ingrediens när man ska göra krukmakeri.
Det verkar som att tjuven bröt sig in genom ett fönster på den övre våningen.
Fienden kastade in nya styrkor i slaget.
Filosofi är inte ett så svårt ämne som du tror.
I klart väder kan vi se ön härifrån.
Plötsligen förlorade kontorsarbetaren sitt temperament.
Du har ett meddelande här.
Den här rörelsen från landbygds- till stadsområden har pågåtts i över tvåhundra år.
Jag föddes och växte upp i landet.
Var snäll och tänd lampan.
Tåget avgick i tid.
Telefonen är trasig.
Kan du kolla om telefonen är trasig?
Oddsen för att Reds vinner är 2 mot 1.
Ge inte upp halvvägs.
Var inte arg.
Det var en tyst natt i vintertid.
De började sälja en ny typ av bil i Tokyo.
Vad är den mest behändliga vägen att ta sig till Tokyo Station?
Det var hans anteckningsbok som blev stulen.
Hur anmäler jag en stöld?
Då hade Tyskland en kraftfull armé.
När jag väl har blivit vald ska jag göra mitt bästa för er alla som har stöttat mig!
Räck upp handen om du vet svaret.
Det var omöjligt att hitta ett svar.
Det var omöjligt att finna ett svar.
Vira en sjal om ditt huvud.
En tiger har rymt från zoot.
En tiger har rymt från djurparken.
Detsamma gäller Japan.
Jag säger samma sak om och om igen.
Ta en karta med dig ifall du skulle gå vilse.
Är du vilse?
Träning är för kroppen, vad läsning är för sinnet.
Det är molnigt.
Molnigt med återkommande regn.
Vilken av de två är tyngst?
Det är en fots längd mellan de två husen.
Jag började tillsammans med två resande kompanjoner.
De två försökte ena efter den andra.
Skär köttet i tunna skivor.
Lägg köttet i kylen, annars kommer det ruttna.
Att föra en dagbok är en bra vana.
Även fast jag satt i solen så kände jag mig kall.
I Japan behöver vi sätta på ett sextiotvåyenfrimärke på ett brev.
Jag är väldigt upptagen hemma.
Vad tycker om Japan?
Vi har många jordbävningar i Japan.
Japans huvudgröda är ris.
Hur många olika pjäser är det i japanskt schack?
Det här är en japansk docka.
Detta är en japansk docka.
En japansk trädgård har vanligtvis en damm.
Japan är varmt och klibbigt om sommaren.
Japan behövde kontakt med västerlandet.
Japan är ett vackert land.
Känner du till någon doktor som kan prata japanska?
Folk säger ofta att japanska är ett svårt språk.
Det finns många amerikaner som kan tala japanska.
Tycker du om japansk mat?
Det är inte alltid lätt att skilja på japaner och kineser.
Vart är den japanska ambassaden?
Efter söndag kommer måndag.
Är det öppet på söndag?
Skulle du vilja spela tennis på söndag?
Vad tycker du om att göra på söndagar?
Vad gillar du att göra på söndagar?
Tålmodighet är den vackraste dygden.
Katten sover på soffan.
Katten sov på bordet.
Katten flydde med en bit fisk från köket.
Brandmannens ansikte var bistert när han kom ut ur det brinnande huset.
Bonde plöjde hans fält hela dagen.
Våg efter våg forsade upp på stranden.
Våg efter våg rullade upp på stranden.
Våg efter våg böljade in på stranden.
Det här är löjligt!
Var inte dum.
Min rygg gör fortfarande ont.
Jag fick en spark i baken.
Du är en ängel som handlar åt mig.
Juryn är oenig.
Är den vit?
Är det vitt?
Explosionen skakade hela byggnaden.
Liftarna var närapå förfrusna när de hittades.
Du passar bra i kort hår.
Boten skall betalas i kontanter.
Brottslingen landsförvisades.
Han är ostoppbar just nu men frågan är hur länge han kan hålla sig kvar vid sin höjdpunkt ut av sin karriär.
Hur lång tid tog det honom att skriva den här romanen?
Detta är hyddan som han levde i.
Jag tycker att det är ganska konstigt att han inte skulle veta någonting sådant.
Vi bryr oss inte om vad han gör.
Det är tydligt att han är hemma.
Han sjöng en sång.
Det är underligt för honom att vara borta från skolan.
Till hans förvåning stannade tåget till kort.
Jag gillar honom.
Hunden följde efter honom vart han än gick.
Jeg vet inte om han kommer att besöka oss nästa söndag.
Vet du varför han skolkade idag?
Vet du anledningen till att han skolkade idag?
Om han hade tagit mina råd så hade han varit rik nu.
Han är säker på att han kommer vinna matchen.
Det tog honom tre månader att lära sig cykla.
Romanerna han skrev är intressanta.
När han log, såg barnen hans långa gråa tänder.
Det är säkert att han kommer att lyckas.
Var är han född och uppvuxen?
Äpplena han skickade mig var utsökta.
Han skickade mig ett föddelsedagskort.
Jag visste att han försökte använda pengarna till att bli guvernör.
Han blir sällan arg.
Jag hade pluggat engelska i två timmar när han kom in.
Ingen vet om han älskar henne eller inte.
Ingen vet vare sig han älskar henne eller inte.
De säger att han har varit död i två år.
Vi vet att han är en modig man.
Vi gör det när han kommer.
Hans försök med att simma över floden misslyckades.
Han misslyckades med att försöka simma över floden.
Hur är han?
Han är min typ!
Om det var han så kunde han gjort sämre ifrån sig.
Det är ingen idé att prata med honom. Han lyssnar aldrig.
Han har god anledning att tro det.
Han verkar förakta folk från Kakogawa.
Han har en bror och två systrar.
Hon har inte mindre än tolv barn.
Han hade tre söner som blev advokater.
Jag borde ha vetat bättre än att ringa honom.
Jag tänkte ringa honom, men jag kom på bättre tankar.
Jag läste brevet åt honom.
Hans stackars hund lever fortfarande.
Hans frånvaro igår berodde på hans förkylning.
Det är knappast värt att bry sig om honom.
Hans skjorta var grå och slipsen gul.
Hans slips matchar bra tillsammans med hans kostym.
Han är längre än sin bror.
Hans dumma svar överraskade allihopa.
Hans dumma svar överraskade alla.
Hans sätt var mycket impopulärt.
Hans otrevliga kommentarer spädde på dispyten.
Hans tal var för kort.
Hans tal fångade vår uppmärksamhet.
Jag tycker inte att hans prestation var något vidare bra.
Hans hus ligger precis över gatan.
Hans hus var litet och gammalt.
Har du hört honom sjunga?
Han uppskattar att det nya huset kommer kosta ungefär trettio miljoner yen.
Han är välavlönad.
Vi trodde att hans hot bara var ett skämt.
Det han sade var inte sant.
Hans fel var avsiktligt.
Hans hobby är att samla på gamla frimärken.
Hans affär orsakade stora förluster.
Hans romaner är för djupa för mig.
Hans bil kolliderade med ett tåg.
Han klär sig som en gentleman, men han talar och uppför sig som en clown.
Hans uppsats är kopplad till min.
Hur stor är han?
Hur gammal är han?
Hans bok blev föremål för kritik.
Hans ilska var förfärlig att se.
Hans uppfinning är överlägsen konventionell utrustning.
Han kände sig obekväm i hans fars närvaro.
Hans rum är alltid i ordning.
Hans svar var kort och koncist.
Hans svar är i princip ett nej.
Jag kan inte stå ut med sin fräckhet.
Hans namn är känt världen över.
Jag hade hans namn på tungan, men jag kunde inte komma ihåg det.
Han var så modig att han inte var rädd för någonting.
Hans historia är sann.
Vi kunde inte godta hans berättelse.
Han berättade inte för John om olyckan.
Han fick sitt vänstra ben skadat i en olycka.
Han har blivit längre och längre.
Han är inte här längre.
Han somnade med radion på.
Även om han säger att han ska återvända till Iran för att gifta sig så är hans planer efter Japan väldigt osäkra.
Han frågade mig vem jag var.
Hans kunskaper i kinesiska gjorde att vi kunde genomföra planen smidigt.
Han är van vid att gå långa sträckor.
Han sa att han hade köpt den boken där dagen innan.
Han går i tionde klass.
Han är tillbaka om tio minuter.
Han tjänar inte mer än femtio dollar i veckan.
Han kommer kunna gå upp och gå om ungefär en vecka.
Han var van att flyga ensam och hade i sin fantasi flugit rutten många gånger.
Han arbetar hårt året runt.
Han är tillbaks om några dagar.
Han bestämde sig inte för att bli författare förrän han var trettio.
Han svarade genom att ge "OK" gesten.
Han såg ut som om han vore sjuk.
Han förstår Er inte.
Han bor i den herrgården.
Det sägs att han är född i Afrika.
Han undersökte Amazonas regnskog.
Han utforskade Amazonas regnskog.
Han genomforskade Amazonas regnskog.
Han är bara en amatör.
Han dricker för mycket.
Han sprang för fort för att vi skulle kunna hinna ikapp.
Jag tror att han är en schyst kille.
Han är från England, men är väldigt dålig på engelska.
Han tog fram några mynt.
Han tog ut några mynt.
Han är alltid full av livskraft.
Han är alltid full av energi.
Han är alltid en man vid full vigör.
Han tappar alltid bort sitt paraply.
Han lämnar alltid sina verk gjorda till hälften.
Han pluggar alltid.
Han studerar alltid.
Han tror fortfarande på hennes ord.
Han gick motvilligt för att träffa henne.
Jag tror att han var arg.
Han gick till affären för att köpa lite apelsiner.
Han rånade en gammal dam.
Han har det bättre än någonsin.
Hans systrar så väl som han själv bor nu i Kyoto.
Han gifte sig med en vacker flicka.
Han har cancer.
Han bestämde sig för att en gång för alla sluta röka.
Han har faktiskt inte ätit kaviar.
Han fyllde glaset med vin.
Han föll aldrig för frestelsen.
Han tycker inte om kaffe.
Han grävde tålmodigt efter fakta.
Han tömde sitt glas.
Han betedde sig som ett barn.
Han har blivit rundare.
Han låter den här pistolen vara laddad.
Han är världens rikaste man.
Han är känd som den bäst advokaten i den här staden.
Han har problem.
Han får komma.
Han spelar golf.
Han fick malaria medan han bodde i djungeln.
Han ådrog sig malaria när han bodde i djungeln.
Jag antar att han kommer tillbaka snart.
Han har redan gått ut.
Hon tycker inte om sport och det gör inte jag heller.
Han hade massor att göra.
Där blev han anfallen av rebellerna.
Han löste korsordet med lätthet.
Han stoppade näsduken i sin ficka.
Han stoppade näsduken i fickan.
Han deltog i mötet.
Han stannade där hela tiden.
Han motsatte sig planen.
Han vårdar de gamla fotografierna.
Han har en stor restaurang nära sjön.
Han skadades allvarligt i trafikolyckan.
Han tog på sig den svarta överrocken.
Han högg ned det där körsbärsträdet.
Han bröt nacken i olyckan.
Han förnekade sin inblandning i historien.
Han beskrev olyckan i detalj.
Han var sen på grund ut av olyckan.
Han förnekade den uppgiften.
Han kunde inte förmå sig att skjuta hjorten.
Han undvek betet.
Han bestämde sig för den röda bilen.
Han skrev ner telefonnumret.
Det tog honom tio minuter att lösa problemet.
Han nämnde det.
Det verkar som att han känner till det.
Han är säker på att det är curry.
Han borde ha varit färdigt nu.
Han verkar inte ha vetat det.
Han håller det hemligt.
Han kunde inte gå längre.
Han vore den sista mannen som skulle göra något sånt.
Han är ofta förskenad till skolan.
Han är ivrig över att tillfredställa allihop.
Han kan ha gått en annan väg hem.
Han har precis kommit hem.
Han är något av en musiker.
Han tycker om att spela tennis.
Han tycker om att se på TV.
Han visste inte vad han skulle göra.
Vart gick han?
Jag tycker inte om honom, för han är slug som en räv.
Han är angelägen att åka dit.
Han pratade väldigt högt.
Han är mycket lång.
Han är mycket lång.
Han var väldigt trött.
Hur länge har han varit borta?
Hur länge har han varit frånvarande?
Han är kortare än Tom.
Han har en Toyota.
Han är duktig med kort.
Han finslipade en kniv.
Han viftade bort flugorna.
Åker han buss till skolan?
Han önskar att han kommer besöka Paris.
Han spelade piano.
Han gick ut trots ösregnet.
Han gör vin av grapefrukt.
Han talar franska.
Han är rädd för ormar.
Han sparkade in bollen i mål.
Han kände i fickan efter tändaren.
Han har skaffat sig vanan att stoppa händerna i fickorna.
Han hade få tänder.
Är han här snart?
Han såg ut som om inget hade hänt.
Han är stolt över att vara musiker.
Har han kommit än?
Han bor inte där längre.
Han har redan gått.
Han är i en desperat sökning efter fler bevis.
Han gjorde äntligen slut med den där kvinnan.
Han är antingen full eller tokig.
Han är bra på rugby.
Han började lära sig spanska genom radion.
Han blåste ut ljuset.
Hon hungrade efter närhet.
Han kände sig fram genom mörkret.
Han är stolt över att vara doktor.
Han är stolt över att vara läkare.
Är han en läkare?
Han är inte en läkare.
Han var själv.
Han var ensam.
Han försökte hårt i förgäves.
Han gör ingenting annat än klagar dagarna i ända.
Han är en slug räv.
Han gick ut i regnet.
Han är en dålig chaufför.
Han är en god simmare.
Han är före i sin engelska klass.
Han stannade upp mitt sitt anförande.
Han var mer än en kung.
Han tycker mycket om musik.
Han gillar musik mycket.
Han tycker mycket om musik.
Han gillar musik mycket.
Vilken tid bad han om ditt svar?
Han har dussintals böcker om Japan.
Han var hemma.
Han promenerade hem.
Han gick hem.
Han är bra på att sjunga.
Han levde inte upp till förväntningarna.
Han har medlemsprivilegier.
Han har gått ut.
Han var inne i sina egna tanker med handen över hans panna.
Han vänjde sig kvickt vid det kalla vädret.
Han vande sig snart vid det kalla vädret.
Av misstag svängde han vänster istället för höger.
Han känner många människor.
Han blev nästan dränkt.
Han var i ett kritiskt tillstånd.
Eftersom han är gift, måste han tänka på framtiden.
Han agerade snabbt och släckte elden.
Han steg på tåget.
Han skyndade sig tillbaka från England.
Han hatar att bli tillsagd att skynda sig.
Han började gråta.
Han krävde att hans lön skulle höjas.
Han har tio kossor.
Han har tio kor.
Han dog i cancer förra året.
Han tycker inte om fisk.
Han bor i Kyoto.
Han är stark.
Han vann matchen tack vare sin starka vilja.
Han ser stark ut.
Han tillgodogjorde det han hade lärt sig.
Han är lärare.
Han längtar efter att bli en lärare.
Han låg på rygg.
Jag råkade höra konversationen.
Han har ett tillräckligt bra omdömde för att inte låna ut pengar till dig.
Han var rädd att du skulle skjuta honom.
Folk säger att han aldrig dör.
Han kommer aldrig att erkänna sin skuld.
Han kommer aldrig att erkänna att det är hans fel.
Han är ogift.
Han blev kry igen.
Han flyttade till en varmare plats med omtanke om sin hälsa.
Han gick ut en runda med hunden.
Han är inte vad han utger sig för.
Han såg en hund i närheten av dörren.
Han räknade ut ljusets hastighet.
Han får göra vad han vill med pengarna.
Han kan göra vad han vill med pengarna.
Han tappade greppet om repet och föll ner i floden.
Han gick inte, och det gjorde inte jag heller.
Han bar sig illa åt.
Han har spelat schack sedan han gick på high school.
Han har ingen stolthet.
Han har en plats i parlamentet.
Vad gör han nu?
Han vill spela fotboll i eftermiddag.
Han satt och läste en bok.
Han skulle aldrig få se sina föräldrar igen.
Han var siste man att komma fram.
Han övertalade sin fru att inte skilja sig.
Han skriver böcker.
Efter att ha misslyckats två gånger i går vill han inte försöka igen.
Han sov gott igårnatt.
Han blev ditsatt för mord.
Han blev falskeligen anklagad för mord.
Han blev snärjd för mord.
Han åker om tre dagar.
Han tabbade sig på jobbet och fick sparken.
Han förnekar ingenting för sina barn.
Han blåste på sina fingrar för att värma dem.
Han kunde lära sig utan instruktioner.
Ska han dö?
Han har en bil som jag gav honom.
Han är lika gammal som jag.
Han önskade att gud skulle välsigna mig.
Han vred om min arm.
Han utövade påtryckningar på mig.
Han lovade mig att vara mer försiktig i framtiden.
Han gav mig ett exempel.
Han visade mig sin frimärkssamling.
Han gjorde mig en trädocka.
Han har gjort sitt yttersta för mig.
Han hittade min cykel.
Han kysste mig på pannan.
Han kollade mig rakt i ansiktet.
Han är min bror, inte min far.
Han stal plånboken av mig.
Han svarade inte på mitt brev.
Han är min chef.
Han beundrade min nya bil.
Han förklarade för min son varför det regnar.
Han är lika lång som min far.
Han behandlar mig som ett barn.
Han känner inte mig.
Han gav oss kläder, och pengar också.
Han är en poet.
Han fuskade under provet genom att kopiera från flickan framför honom.
Han kommer inte att misslyckas vid examinationen.
Han är inte för fattig för att köpa en cykel.
Han kopplade på husvagnen på sin bil.
Han sökte i sin väska efter bilnyckeln.
Där såg han det han hade drömt om.
Han stack sitt hus i brand.
Han satte eld på sitt hus.
Han jobbade hårt för att försörja sin familj.
Han är medveten om hans eget fel.
Han erkände sina misstag.
Han skrev ner sina tankar i sin anteckningsbok.
Han ägnade all sin tid till att studera historia.
Han väntade på sin tur.
Han kan inte ens skriva sitt eget namn.
Han trodde inte sina ögon.
Han förklarade hans situation för mig.
Han förklarade sin situation för mig.
Han tog sig friheten att skriva till damen.
Han har ett bra rykte som affärsman.
Han förklarade varför experimentet misslyckades.
Han är social av sig.
Han tvättar bilen.
Han har sålt sin bil, så han tar tåget till kontoret.
Han verkar ha haft ett svårt liv i sin ungdom.
Han ser ung ut.
Han lider av en svår sjukdom.
Han stannade hos hans fasters hus
Han stannade hos hans mosters hus.
Han sov över hos hans fasters hus.
Han sov över hos hans mosters hus.
Han förklädde sig till en kvinna.
Han gifte sig med en skådespelerska.
Han tillverkade en liten hundkoja.
Han siktade mot fågeln.
Han ser lite trött ut.
Han kallades att vittna.
Han brände hål i rocken.
Han kom till New York för att söka jobb.
Han arbetar fortfarande i arbetsrummet.
Han är nöjd med sin nya bil.
Han berättade sanningen.
Han sade sanningen.
Han är en gentleman.
Han verkar snäll.
Han är medveten om faran.
Han gillar skvaller.
Han är oerhört stilig.
Han klarade det.
Han hann.
Han är av naturen en vänlig person och populär hos barnen i området.
Han sa åt eleverna att vara tysta.
Han ägnade sig helt helhjärtat åt henne.
Han var inte samma glada man han en gång var.
Han blev tilldelad en ansvarsfull position.
Är han en lärare?
Han drunknade i floden.
Han bor på andra sidan floden.
Han gick inte upp tidigt.
Han steg inte upp tidigt.
Han är sitt vanliga jag.
Hon började springa.
Han höll andan.
Han måste köpa en ny cykel åt hans son.
Han var så upptagen att han skickade sin son istället för att gå själv.
Han är grov till sättet.
Han befordrades till överste.
Han är en storätare.
Han valdes till president.
Han greps för skattefusk.
Jag såg på honom att han bara låtsades läsa.
Han har skrivit en bok om Kina.
Han tror på det övernaturliga.
Han rensade gatan på kastanjer.
Han tjänstgjorde utan allvarligare anmärkningar till han uppnådde pension.
Han studerar astronomi, eller stjärnlära.
Han längtar efter stadsliv.
Han ansträngde sig ej.
Han är stolt över att ha tagit examen vid Tokyo Universitet.
Han var intresserad av Orientens mysterium.
Hans huvud värkte.
Han måste komma söderifrån.
Han har setts som Japans svar på Picasso.
Han vet bättre än att gifta sig med henne.
Han är bra på att imitera hennes irländska brytning.
Han tog henne i handen.
Han höll henne i ärmen.
Han tog med henne till vårt ställe.
Han ser trött ut.
Verkar som om han är trött.
Han verkar trött.
Det verkar som att han är trött.
Han blödde näsblod.
Han kunde inte komma tillbaka, då han var sjuk.
Han har tre familjemedlemmar att försörja.
Han är bara en vanlig kontorsråtta.
Han står på scenen.
Han tvingade sig in i rummet.
Han rusade in i rummet.
Han hade en underlig dröm.
Han kommer att gå.
Han behöll hatten på.
Han var upptagen.
Han var arg över att jag hade kränkt honom.
Han frågade mig om jag ville åka utomlands.
Han lämnade boken på bordet.
Han skulle hellre dö än att gå upp tidigt varje morgon.
Han åker skidor i Hokkaido varje vinter.
Jag somnade.
Han är en man att räkna med.
Han är en man som man kan räkna med.
De förklarade sig oskyldiga.
Han använde hennes cykel utan att fråga om lov.
Han kysste sin dotter på pannan.
Han högg av en gren från trädet.
Han blev blind.
Han satt där med sina ögon stängda.
Han är galen i baseboll.
Han är väldigt upptagen med att skriva till hans vänner.
Han drog förbi en vän.
Han blev en berömd sångare.
Han drog sig tillbaks till sitt rum efter kvällsmaten.
Han visste inte vad han skulle göra med den överblivna maten.
Han kommer att komma.
Han är på väg och kommer att anlända i sinom tid.
Han bor med sin föräldrar.
Han skrev till sina föräldrar.
Han klagade över att rätten smakade dåligt.
Han utförde arbetet så gott han förmådde.
Han sprang inte tillräckligt fort nog för att hinna med tåget.
Han talade inte såvida han inte blivit tilltalad.
Han erkände att han hade tagit mutor.
Han lever i lyx.
Vi visste inte vilket tåg de skulle vara på.
Jag bryr mig inte om vad de säger.
De har ingen annanstans att gå.
De har ingen annanstans att ta vägen.
Ett slagsmål började utan någon anledning mellan dem.
De skillde sig förra året.
Deras trädgård är full ut av väldigt vackra blommor året runt.
Deras nationalism var en ut av orsakerna till kriget.
De dricker coca-cola.
De är skådespelare.
De är korta och smala.
De är korta och smala.
De har tolv barn.
De lyssnar inte alltid på sina föräldrar.
De lyder inte alltid sina föräldrar.
Nu har de tre barn.
De bor i en liten by i England.
De erbjöd gästerna lite kaffe.
De frågade Kate om hon kunde sitta barnvakt åt barnet.
De döpte hunden till Shiro.
De såg efter pojken.
De kommer att komma överens på den punkten.
De hatade Tom.
De stod på rad.
De erbjöd assistans.
De erbjöd hjälp.
De är ivriga på att få veta vad som hände.
De är spända på att få veta vad som hände.
De har alla självständiga betydelser.
De har en gemensam hobby.
De passar varandra på grund ut av deras närliggande intressen.
De bestämde sig för att bygga en bro.
De byggde en bro.
De bor i ett nytt hus nära parken.
De är gymnasieelever.
De plaskade vatten i mitt ansikte.
De lät mig vänta länge.
De har något gemensamt.
De gick hand i hand.
Skriver de ett brev?
De kämpade för religionsfrihet.
De är nöjda med det nya huset.
De tackade Gud.
De skymtade mannen genom folkmassan.
De leker gärna i snön.
De är lärare.
De seglade runt världen.
De försökte fly.
De gratulerade honom till hans bröllop.
De gjorde honom till klubbens ordförande.
De ser honom som en hjälte.
De togs till fånga.
De är lika starka som vi.
De skrattade åt min idé.
De kommer inte förrän imorgon.
De gifter sig nästa månad.
De kan tänka och tala.
Låt honom vänta ett ögonblick.
Låt honom vänta ett slag.
Jag måste hjälpa honom.
Jag vinkade av honom vid flygplatsen.
Det är dumt av dig att tro på honom.
Känner jag honom?
Det går inte att förväxla honom med hans lillebror.
Hon kan prata tio språk.
Hon köpte en bok i affären.
Precis när hon skulle lämna affären så såg hon en vacker klänning i fönstret.
Jag var irriterad över att hon fortfarande sov.
Har du hört av henne?
Det är dig som hon älskar, inte mig.
Fråga henne vad hon har köpt.
Jag fick reda på var hon var.
Mannen som hon ska gifta sig med är en astronaut.
Jag tog det förgivet att hon skulle hålla med mig.
Hon kan bara lita på honom.
Jag lade märke till att hon satt på främsta raden.
Jag lade märke till att hon satt på första raden.
Vem hon är har jag ingen aning om.
Inte underligt att hon inte dök upp för att ge honom ett avsked. De har gjort slut.
Det är inte för att hon är vacker som jag gillar henne.
Det slog honom aldrig att hon skulle bli arg.
Ge henne det här brevet när hon kommer.
Var såg du henne?
Trots alla hennes brister gillar jag henne.
Skall du presentera mig för henne?
Var snäll mot henne.
Var snäll mot henne, Bill.
Hennes far avled i förra veckan.
Jag känner henne inte alls.
Hennes klänning såg billig ut.
Hennes engelska är utmärkt.
Hennes ansikte blev rött plötsligen.
Hennes argument byggde inte på fakta.
Hennes ledighetsansökan avslogs.
Hennes storasyster gifte sig förra månaden.
Nyheten om hennes död kom som en blixt från klar himmel.
Hennes skämt gick inte hem.
Hennes röst går mig på nerverna.
Min mormor blev åttioåtta år gammal.
Jag kan inte ta hennes plats som engelsklärare.
Hennes hår är långt och vackert.
Färgen av hennes klänning och skor matchade varandra bra.
Hennes namn är känt världen över.
Tårar föll från hennes ögon.
Hennes enda fritidsintresse är att samla på frimärken.
Hennes enda önskan var att träffa sin son igen.
Hon är en kontorskvinna.
Hon tycker om vin.
Hon gillar vin.
Hon dog 1960.
Hon kom inte innan två.
Hon kom inte förrän två.
Hon spelade piano tillräckligt bra.
Hon höll just på att skära upp gurkor.
Hon behöver hjälp.
Hon var försiktig med att inte slå sönder glasen.
Hon kan spela den här melodin på piano.
Hon föll ner för stegen.
Hon fortsatte prata.
Hon ville gifta sig omedelbart.
Hon har blivit en helt annan person.
Hon rörde om i kaffet med en sked.
Hon valde skorna som passar till klänningen.
Hon valde skorna som matchar klänningen.
Hon betalade sju procents ränta på lånet.
Hon frågade var huset låg.
Hon började prata med hunden.
Hon blev väldigt arg på barnen.
Tanken på att hon skulle möta den berömda sångaren fick henne att rysa av spänning.
Hon sa att hon inte gillade den, men jag tyckte, personligen, att den var väldigt bra.
Hon översatte det ord för ord.
Hon slöt in det i papper.
Hon har en del egna pengar.
Hon har äntligen nått Arktis.
Hon äter middag nu.
Hon tillhör tennisklubben.
Hon älskar att se på tennismatcher på TV.
Jag undrar varför hon inte berättade om det för honom.
Överallt hon kommer är hon uppskattad.
Hon är mycket vacker.
Hon älskar Tom.
Hon gråter.
Hon är långt ifrån dum.
Hon log.
Hon hade hjärtformade örhängen.
Hon räckte upp handen för att få bussen att stanna.
Hon talar tillräckligt tydligt för att vara lätt att förstå.
Hon skrek i sin förvåning.
Hon skrek till av förvåning.
Hon valde ut en rosa skjorta för mig att prova.
Hon erkände att hon inte kunde prata franska.
Kan hon franska?
Talar hon franska?
Hon gillar klassiska kompositörer såsom Beethoven och Bach.
Hon är väldigt rädd för ormar.
Hon är min flickvän.
Hon har inte kommit hit än.
Det dröjer inte länge innan hon är tillbaka.
Hon pratar om Paris som om hon har varit där flera gånger.
Hon pratar engelska som om det vore hennes modersmål.
Hon går sällan ut.
Hon försökte hoppa upp en andra gång.
Hon är ute efter ett bättre jobb.
Hon är sig själv igen.
Hon var tvungen att ge upp planen.
Hon hade en radio.
Hon kom ensam.
Hon är för ung för att skaffa körkort.
Hon är en god simmare.
Hon kan inte bara prata engelska utan också franska.
Hon kan inte bara tala engelska, utan också franska.
Hon kan prata både engelska och tyska.
Hon studerade utomlands för att borsta upp hennes engelska.
Vad har hon?
Hon talar inte japanska hemma.
Hon pratar inte japanska hemma.
Är hon hemma?
Hon gick hem.
Hon har satt sitt hus till försäljning.
Hon sjunger bra.
Hon gillar att prata framför oss.
Hon instämmde med våra begär.
Hon har en stuga vid havet.
Hon skyndade ner för trapporna.
Hon är inte så ung som hon ser ut.
Hon är pigg på att sticka utomlands.
Hon gick ut.
Hon rynkade pannan.
Hon är en sjuksköterska.
Hon är inte sjuksköterska, utan läkare.
Hon verkade inte intresserad.
Hon var nära på att drunkna.
Hon är utom sig av glädje.
Det verkade som om hon redan hade fått pengarna.
Hon går ofta och shoppar på helger.
Hon betalade för att gå på konserten.
Hon såg upp mot himlen.
Hon är lika lång som du.
Visade hon dig bilden?
Hon är på intet vis självisk.
Är hon gift?
Hon är inte gift.
Hon är fem år gammal.
Hon är lycklig.
Hon beställde en kopp te.
Hon var klädd i svart.
Hon böjde sig ner.
Hon var på vippen att gråta.
Hon var gråtfärdig.
Hon var gråtfärdig.
Hon var på väg att svimma.
Hon såg mer vacker ut än någonsin förrut.
Hon är ute nu.
Jag har en känsla på mig att hon kommer att komma idag.
Hon satt och rökte.
Hon kom sist.
Medicinen var hennes sista utväg.
Igår hon köpte grönsaker.
Hon lämnade scenen förra året.
Hon var på humör för en promenad.
Hon har en viktig roll i vår organisation.
Hon kanske berättade en lögn för mig.
Hon gav mig de här gamla mynten.
Hon meddelade mig om hennes avfärd.
Hon frågade mig om jag mådde bra.
Hon är min typ.
Hon nekade mitt önskemål.
Hon känner mig.
Hon undviker mig.
Hon har en väldigt prydlig handstil.
Hon kommer aldrig i tid.
Hon fick en stor summa pengar i förskott för hennes nästa roman.
Hon övergav sina barn.
Hon kände sig illa till mods vid tanken på hennes framtid.
Hon skämdes för sin obetänksamhet.
Hon är stolt över sin dotter.
Hon brann med svartsjuka.
Hon har en bild.
Du borde ha bett om ursäkt till henne.
Hon måste ha varit väldigt vacker när hon var ung.
Hon borde ha gjort klart sina läxor.
Hon kan vare sig läsa eller skriva.
Hon ser sin chef som sin far.
Hon är mörkhyad.
Hon har gått och lagt sig.
Hon valde en hatt som matchade hennes klänning.
Hon är snäll.
Hon var snäll och tog mig till sjukhuset.
Hon är tystlåten.
Hon är tyst.
Hon bar babyn på ryggen.
Hon är väldigt duktig på att imitera sin lärare.
Hon är tvilling.
Hon ger sin son för mycket pengar.
Hon köpte en kamera till sin son.
Hon klappade sin son på axeln.
Hon har tagit på sig alltför mycket arbete.
Hon vann första pris i en matätartävling.
Hon svor högt.
Vem är hon?
Hon blev arg.
Hon gick ut.
Hon ser ung ut för sin ålder.
Hon läste hans brev om och om igen.
Det hade aldrig slagit henne att han skulle bli bestraffad.
Hon ser fram emot att få träffa honom igen.
Hon sa att de var goda vänner till henne.
Hon ville hjälpa dem.
Hon vill hålla honom på avstånd.
Hon måste hjälpa honom.
Hon ser ledsen ut.
Hon såg ledsen ut.
Hon har en fin docka.
Hon kunde inte komma för hon var sjuk.
Fattig som hon var gav hon honom det lilla hon hade ut av sina pengar.
Hon var på dåligt humör.
Hon lever ett olyckligt liv.
Hon hjälpte sin far med trädgårdsarbetet.
Han ska övertala sin far att köpa en ny bil.
Hon har sönder något varje gång hon städar rummet.
Hon sa att hon hade en förkylning.
Hon kunde inte hindra sin dotter från att gå ut.
Hon gav mig inte sitt namn.
Hon kom in helt tårögd.
Hon lever på grönsaker och råris.
Hon var modig.
Hon blir sen till maten.
Hon kanske inte kommer.
Kommer hon att komma?
Hon är mer vis än smart.
Hon antydde att hon kanske skulle studera utomlands.
Hon bad mig att se efter hennes bebis medans hon var borta.
Hon såg till att resenären hade mat och kläder.
Hún eldar illa.
Hon bytte ämnet.
Hennes arm är gipsad.
Kommer hon med?
När såg du henne senast?
Känner du henne?
Han kramade henne.
De tittade på teve.
De tittade på tv.
De vann faktiskt.
De stack vid klockan 5, så de borde vara hemma vid 6.
Du ser sjuk ut.
Till hennes sorg hade hennes son lämnat henne ensam.
Var inte ledsen.
Är du trött?
Kan du hålla det en hemlighet?
Jag såg ett flygplan.
Har du redan bokat våra platser på flygplanet?
Flygplan kan höras långt före de syns.
Min näsa kliar.
Prinsessan låg och blundade.
Isen smälter.
En sjukdom förhindrade honom från att gå ut.
Fast han är mycket fattig, är han ändå för god för att ljuga.
Tyvärr gick guiden fel.
Det är allt annat än omöjligt.
Det är inte lönt att klaga.
En dam, vars man är en känd forskare, kom över från den andra sidan.
En kvinna vars man har dött är en änka.
Var ligger damernas?
Kom så skakar vi mattan.
Vart gick pappa?
Min fars bil är gjord i Italien.
Min far hade redan varit en gång i Grekland.
Min far röker.
Min far lagade en trasig stol.
Min pappa insisterade på att vi skulle vänta på tåget.
Min far insisterade på att vi skulle vänta på tåget.
Min far är inte hemma.
Min far besökte min farbror på sjukhuset.
Min far älskar min mor.
Det besegrade laget lämnade så sakta planen.
De sårade kom med ambulans.
Det var många människor i rummet.
De smyckrade upp rummet med blommor.
Du måste städa ditt rum.
Jag skulle vilja byta rum.
Vinden blåste hela dagen.
Var försiktig så att du inte blir förkyld.
Har den ett badrum?
Tog du ett bad?
Jag gav det ett försök och tänkte att allting är värt ett försök. Men att sätta ihop ett sånt här program har jag ingen chans för.
Man måste dra gränsen någonstans.
Fysik är mitt favoritämne.
Jag vet.
Meningar börjar med en stor bokstav.
Sluta klaga och gör som du blivit tillsagd.
Lyssna på detta!
Vet du vad?
Det fanns en hatt och en kappa på vägen.
Du behöver inte vara rädd. Han kommer inte att göra dig illa.
Ge mig ett exempel till.
Visa mig ett annat exempel.
Det är konstigt.
Jag hör ett konstigt ljud.
Jag vill ha pengarna tillbaka.
Prata med mig!
Avdokaten insisterade över klientens oskyldighet.
Advokaten förklarade den nya lagen för oss.
Min mor är ute.
Mor går till sjukhuset på morgonen.
Mamma var allt som oftast väldigt upptagen.
Mor, far. Titta på ert lilla monster.
Mor köpte två flaskor apelsinjuice.
Hjälp mig lyfta paketet.
Många barn stannar efter skolan för klubbaktiviteter.
Min hat trillade av.
Häng din hatt på kroken.
Glöm inte att signera med ditt namn.
Glöm inte att skriva under med ditt namn.
Han skrev ner det för att inte glömma det.
Man har funnit olja under Nordsjön.
Jag betalar notan.
Jag har rätt.
Vi spelade schack inte så mycket för att vi gillade att spela som för att bara slå ihjäl tiden.
Min lägenhet är i närheten.
Min lägenhet ligger här i närheten.
Förstår du vad jag menar?
Min far är så att säga en vandrande ordbok.
Jag är inte trött alls.
Jag gillar jazz.
Jag är så lycklig.
Jag har aldrig ätit mango förut.
Jag kan inte vänta längre.
Jag måste bege mig nu.
Jag måste gå nu.
Jag måste bege mig nu.
Jag är trött på att äta på restaurang.
Jag är i London.
Jag är vänsterhänt.
Jag har två bilar.
Jag är ung.
Som pojke brukade jag ligga på gräset och titta på de vita molnen.
Jag vill sova.
Jag växte upp på landet.
Jag är förkyld.
Jag också.
När kan vi äta?
Jag har inte tid att läsa.
Är det sant?
Det känns som att jag är på bättringsvägen.
Om jag visste sanningen skulle jag ha berättat den för dig.
Hur är det med din syster?
Min syster leker med dockan.
De hämtar våra sopor varje måndag.
Att träna varje dag är nödvändig för din hälsa.
Jag tycker inte om att handla varje dag men jag måste göra det.
Kan jag få en kudde?
En av fördelarna med att bo i en demokrati är att man får säga vad man tycker och tänker.
Jag kunde inte sova.
Är det gratis?
Reta inte honom bara för att han inte kan skriva sitt namn.
Det är inte den typen av sjukdom som sätter ditt liv i fara.
Akiko har några vänner i Frankrike.
Jag ska fråga honom om det imorgon.
Jag ska ringa om det imorgon.
Vädret ska bli bättre imorgon.
Jag tror inte att det kommer att regna i morgon.
Det är söndag imorgon.
I morgon ska jag gå och shoppa.
Imorgon är det hennes föddelsedag.
Imorgon fyller hon år.
Vi ska ha prov i engelska imorgon.
Vi ses i skolan imorgon.
Bomull absorberar vatten.
Det är intressant.
Det är rea på pälskappor.
Kan du ge mig en filt?
För träd är grenar vad lemmar är för oss.
Löven virvlade runt i gården.
Kimura joggade i parken varje dag.
Håll käften, eller så slår jag ner dig.
Mina ögon är ömma.
Jag är vaken.
Blunda och sov.
Komm tillbaka!
Poängen är huruvida hon kommer att läsa brevet eller ej.
Är det utegångsförbud?
Dagen gryr.
Det var natt.
Det är roligt att spela baseball.
Jag vill att du håller ditt löfte.
Är du allergisk mot någon medicin?
Förklara hur man tar medicinen är du snäll.
Kastrullen kokar.
Han är snäll.
Till och med en bra dator kan inte klå dig på schack.
Jag sov inte igårnatt.
Det är middagsdags.
Jag behöver en extra kudde.
Finns det reserverade platser på tåget?
Den misstänkte ljög för polisassistenten.
Du kan komma med oss om du vill.
Snälla kom.
Kom snälla du, jag är ivrig över att se dig.
Kom och hjälp oss.
Håll utkik efter hans senaste film som kommer ut nästa månad.
Jag skulle vilja träffa dig igen nästa vecka.
Memorera dikten till nästa vecka.
Det går inte att förutsäga vad som kommer hända nästa år.
Jag kommer att kunna träffa honom nästa år.
Hästens fall resulterade i ett brutet ben.
Koka ett ägg.
Det är lättare att lyfta än att landa.
Stå upp.
Ställ dig inte upp.
Kan du ta hand om våra husdjur medan vi är borta?
Kan ni ta hand om våra husdjur medan vi är borta?
Har du badat än, Takashi?
Nöjet av att resa runt är vanligt hos nästan alla personer.
Nyheten om de två företagens sammanslagning kom ut igår.
Båda föräldrarna lever fortfarande.
Det var svalt och skönt, men nu börjar det bli kallt.
Kan jag få ett kvitto, tack?
Midori åt flest apelsiner.
Pojken som bor här intill kommer ofta hem sent.
Vem är det som bor här intill?
Grannhunden skäller alltid.
När hennes grannar var sjuka frågade hon doktorerna att ge dem medicinska hjälpmedel.
Vi besökte historiskt intressanta platser.
Tåget avgår om tio minuter.
Vi hinner med tåget.
Tåget var fullt med passagerare.
Tåget försenades av snön.
Kärlek och hosta kan inte döljas.
Kärleken är till sin natur blind.
Tack för att du tog mig hit.
Hör av dig!
Den gamle mannen och Sjön är en väldigt spännande bok.
Det är en självklarhet att grundläggande mänskliga rättigheter bör respekteras.
Har du någonsin ätit japansk mat?
Prata inte!
Jag svettades under armarna.
Bränt barn skyr elden.
Man ska inte väcka en sovande orm.
"Om det är pengar så lånar jag inte ut något" sa jag kort och gott.
Ah, är det så att du blir generad över att bli kallad vid ditt första namn?
Han inser inte att han är tondöv.
Bortsett från hans häl så var Akilles odödlig.
Det beror på, förstår du, att jag har vetat sen länge att han inte är den sortens människa.
De här reporna syns väldigt mycket så jag skulle vilja få dom reparerade.
Tack vare Harunas "väder läge" blev Kaoris iver väldigt dämpad.
Pandor bor i bambusnår.
Helens ord fyllde mig plötsligt med ny energi.
Helens ord fyllde mig plötsligt med ny kraft.
När jag frågade honom efteråt verkade det som han inte hade menat det som ett skämt.
På grund av några oundvikliga omständigheter i sommar kan jag inte bo i min semesterstuga.
Till och med under arbetstid ger jag i lönndom efter för mitt internetberoende.
Hur sent kan jag ringa?
Att förlora min dotter har berövat mig livsglädjen.
Han har kommit att se ut att vara en rävaktig premiärminister som utnyttjar makten i sitt ämbete till fullo för egen vinning.
Alle man, överge skeppet!
Hela besättningen, överge skeppet!
I svåra sorgfyllda tider, låt oss då göra något för andra.
Det nuvarande lösenordet är "eosdigital".
Av någon anledning fungerade inte mikrofonen tidigare.
Om du strular till det så kan det inte göras om, så strula inte till det!
Jag har problem med att pulvermedicin.
Dock är det något som överlevandena inte känner till.
Förlåt, jag hade inte med det att göra.
Hela familjen hjälpte till med att skörda vetet.
Då är det dags för din halshuggning. Har du inga sista ord?
Min son som går i femteklass har förflyttat sig till skolan i Nagoya från Shizuoka.
Vilket land kommer du ifrån?
Jag vill köra ett Windows 95 spel.
Kan du förklara hur diskmaskinen fungerar?
Han är lika gammal som jag.
Om det är gratis, ta så mycket du kan.
Jag borde sluta skjuta upp saker och ting.
Jag är kines.
Kaffe och cigaretter.
Jag har sett en artikel på Tatoebabloggen om en ny version som ska komma ut snart. Har du läst den?
Kan du hjälpa mig att översätta dessa meningar till kinesiska?
Du kan inte döda dig själv genom att hålla andan.
Vem är han?
Lite tidigare imorse fick jag ett enanstående nådigt samtal från senator McCain. Senator McCain kämpade länge och hårt i den här kampanjen. Och han har kämpat ännu längre och hårdare för det land han älskar. Han har stått ut med uppoffringar för Amerika som de flesta av oss inte kan föreställa sig. Det vore bättre om vi var i tjänst framställd ut av denna modiga och osjälviska ledare.
Jag är inte på väg någonstans.
Jag är gravid.
Jag vet inte.
När man är i Rom så gör som romarna gör.
Ta seden dit man kommer.
De är alla oskyldiga barn.
Studera de här meningarna.
Vi singlar slant om det.
Han förstod inte hennes skämt.
Vem är du?
Det var bara ett skämt.
Den såg billig ut.
Det såg billigt ut.
Vi ses!
Hej då.
Gott Nytt År!
Jag spelar fiol.
Jag är vegetarian.
Jag äter inte kött, fisk, skaldjur, fjäderfän eller buljong.
Dörren är öppen.
Gick du i skolan idag?
Jag älskar arabiska.
Varifrån kommer du?
Var är ditt hus?
Var bor du?
De är mina bröder.
Bilal är utbildad.
Är du lärare eller student?
Han är sjuk.
Jag kommer från Norge.
Vet du om han kommer till festen?
Har du skrivit upp telefonnumret?
Har du skrivit ned telefonnumret?
Solen skiner.
Den här boken verkar intressant.
Denna bok verkar intressant.
Den här boken handlar om Kina.
Eleverna lyssnar på en historieföreläsning.
Katter tycker inte om vatten.
Jag pratar inte tyska.
Det är hett idag.
Det är hett idag.
Förlåååt. Jag kunde inte sova i går kväll, så jag försov mig. Hihi!
Vi ska se.
Hej.
Jag var försenad på grund av trafiken.
Tack!
Vad gjorde du?
Såg du blicken han gav mig?
Hans mål är att bli en lärare.
Städa rummet.
Jag är högerhänt.
Latin är ett dött språk.
Prata inte strunt.
Jag måste lämna dig.
Jag kommer inte ihåg ditt namn.
Du känner dig ensam, eller hur?
Vi har tre flygplan.
Datorn är en komplicerad maskin.
Det är lite kallt idag.
Han torkade svetten från ansiktet.
Jag känner henne inte.
Han är lång och stilig.
Hon hatade honom.
På bussar bör ungdomar ge sina sittplatser till de äldre människorna.
Hon ringde mig flera gånger.
Hon blev påkörd av en bil.
Hon kommer kanske.
Mary kom in.
Han ljög för oss.
Han tycker om att se på TV.
Det är bara ett par få minuter kvar tills tåget går och hon har inte dykt upp än!
Vi är män.
Kanske förstår hon senare vad jag menade.
Jämfört med hans far är han väldigt ytlig.
Alla säger att han ser ut precis som sin far.
Jag har bestämmt mig för att vara glad för det är bra för min hälsa.
Han älskar att resa.
Jag känner på mig att han känner till hemligheten.
Jag förstod inte hans skämt.
Vad är detta?
Jag har inte hört något från honom sen dess.
Sömnbrist är inte bra för kroppen.
Det är omöjligt att inte bli fascinerad ut av hans skönhet.
Jag ska gå rakt på sak. Du får sparken.
Alla djur är lika, men vissa djur är mer lika än andra.
Enligt tidningen begick han självmord.
Sommaren är över.
Han älskar henne.
Jag träffade just henne på gatan.
Jag träffade henne på vägen till skolan.
Jag känner mig inte för att träffa henne nu.
Vad är det för skillnad mellan en by och en stad?
Ju mer du lär känna henne, desto mer kommer du att gilla henne.
Giraffer har mycket långa halsar.
Det var lätt att hitta hans kontor.
Du verkar frånvarande.
Vill du gifta dig först eller skaffa barn först?
De är alla kannibaler här, utom mig, jag bara blir uppäten.
Jag cyklade enhjuling idag.
Det här är hans bil, tror jag.
Detta är hans bil, tror jag.
Har du ett recept?
Tack!
Tack!
Tack!
När jag tänker på de där eleverna får jag huvudverk.
Hej världen!
Jag går alltid.
Jag kom från Kina.
Hon tycker om rysk pop.
Jag tror inte att han kommer.
Han är smart.
Han är intelligent.
Jag lade på och ringde henne igen.
Jag vill tillbaka nu.
Vi kunde inte gå ut på grund av tyfonen.
Vad vill du dricka?
Vad skulle du vilja äta?
Vilken föredrar du? Den här eller den där?
Vi stötte på dem vid bussterminalen.
Vår engelsklärare är både sträng och snäll.
Min engelska är inte alls bra.
Han blev polis.
Det finns få webbsidor på tatariska på internet.
Nästa koncert kommer att hållas i Juni.
Jag kommer så fort jag kan.
Far, får får får? Nej, får får lamm.
Tomten stod på tomten
Vad gjorde du i går kväll?
Vad gjorde du i helgen?
Vad gjorde du i går kväll?
Under den stalinistiska eran blev fångar i koncentrationsläger slavar i statens tjänst.
Enligt väderprognosen ska det snöa i morgon.
När lämnar din far hans kontor?
Vad äter vi ikväll?
Strax innan bröllopet skrek den berusade fadern: "Jag kommer inte att lämna ut min dotter till någon främling!" till brudgummen.
Enligt många religioner är äktenskapsbrott ett brott.
Det är inte en fru jag vill ha, utan en knullkompis.
Jag tycker om att gå och titta på baseboll.
Förstår du mig?
Var är flygplatsen?
Var ligger flygplatsen?
Var snäll och tala långsamt.
Är mjölken god?
Vilken tand gör ont?
Borde jag köpa någonting till honom?
Grekerna äter också ofta fisk.
Hur länge kommer du att vara i Japan?
Du är den sista personen jag förväntade mig att träffa här.
Vad hände på bussen?
Många tror att jag är tokig.
Stäng dörren.
Market Square är det historiska centret i staden.
Som man bäddar, får man ligga.
Tom är en bra person
Det kommer antagligen att snöa i morgon.
Det här året erbjuder vi samma språkkurs som i fjol.
Mitt språk är inte med på listan!
Vad heter du?
Vad är ditt namn?
De säger att han föddes i Tyskland.
Det sägs att han föddes i Tyskland.
Jag är hungrig.
Jag är hungrig.
Jag är bäst.
Jag är bäst.
Vad skulle världen vara utan kvinnor?
Du måste vara på stationen senast klockan fem.
En gång fann jag en bok där.
Du kan lita på honom.
Vilket tåg tänker du ta?
Jag har en katt och en hund. Katten är svart och hunden är vit.
Gör som du vill.
Har jag fel?
En man kan leva och vara frisk utan att döda djur för mat. Därför deltar han i att ta djurs liv enbart på grund ut av hans aptit om han äter kött, och att bete sig så är omoraliskt.
Det viktiga är inte hur en man dör, utan hur han lever.
Säg mig vad du äter, så ska jag säga dig vad du är.
Jag betalar.
Varför var du där?
Jag bad henne att vänta ett slag.
Vi får se vad som händer.
Deras kontor visade sig ha många kvinnor.
Ann gillar choklad.
Ann tycker om choklad.
Det är okej.
Var snäll och kom och hjälp mig.
Vad är detta?
Var snäll och sätt på dig skorna.
Provresultatet visade hur mycket han hade pluggat.
Sten, sax, påse.
Varsågod och sitt ner.
Jag har inga pengar.
Allt i denna värld är blott en dröm.
Han blev av med sitt jobb.
Mina ögon gör ont.
Jag läste just ut Svindlande höjder.
Två personer kommer in på den här biljetten.
Vi har mycket snö vintertid.
När kommer ni att gifta er?
"Hur gammal är du?" "Jag är sexton år."
För länge sedan fanns det en bro här.
Tv:n är på.
Jag skulle vilja ha något att dricka.
Jag började att läsa boken.
Alister dödade Barbare.
Mary hjälpte sin mor att laga mat.
Mary hjälpte sin mamma att laga mat.
Betty är danslärare.
Hur kan folk sova på planet?
Hur lyckas folk sova på planet?
Vi spelar ofta schack.
Det enda gången då folk inte tycker om skvaller är när du skvallrar om någonting om dem.
Vänta, skojar du? Varför skulle vi vilja åka till en sådan avlägsen plats?
Dubbelklicka på ikonen.
De fångade rävar med fällor.
Han var i Frankrike.
Vad vet du om honom?
Schweiz är ett väldigt vackert land och är mycket värt att besöka.
Han är amerikan ut i fingerspetsarna.
Han vände bort blicken.
Jag använder Firefox.
Jag är ledsen, vi har helt slut på manti.
Jag var lärare.
Om du vill ha fred, förbered dig för krig.
Jag förstår.
Det stämmer!
Gå iväg.
Självklart.
Ursäkta mig.
Det är mitt jobb.
Säg det tydligt.
Försök en gång till.
Jag är mänsklig.
Jag är människa.
Jag är en människa.
Jag har ingen pengar.
Titta bakom dig.
Det är en fin dag.
Detta är ett litet steg för en människa men ett jättekliv för mänskligheten.
Jag är seriös.
Det är lunchdags.
Kom med oss.
Självklart!
Jag mår bra.
Jag är mätt.
Jag är väldigt upptagen.
Ett kuvert och ett frimärke, tack.
Är du hungrig?
Är ni hungriga?
Vilken skitstövel!
Behöver jag någon medicin?
Behöver jag opereras?
Sysslar du med någon sport?
Har du barn?
Har du skor och strumpor?
Kommer du ihåg oss?
Kasta ingenting på marken.
För Guds skull.
Knulla din mamma.
Har posten kommit än?
Han är arton månader gammal.
Han är en av Spaniens mest kända författare.
Han tycker om att simma.
Han behöver en stege.
Han kastade ut mig ur huset.
Hjälp!
Den är för stor.
Länge leve Sovjetunionen!
Lugna ner dig.
Lugna ner er.
Han kan också tala ryska.
Du måste inte äta.
Livet är roligt.
Städa ditt rum.
Det är gratis.
Jag har blivit bättre.
Hur vet du det?
Vad kostar en öl?
Hur gammal är du?
Hur gammal är din son?
Hur stavar man ditt efternamn?
Hur stavar man ert efternamn?
Jag är Lin.
Jag är inte intresserad.
Jag har ryggont.
Jag har ont i ryggen.
Jag behöver ett jobb.
Jag behöver en anteckningsbok för att föra mina anteckningar.
Jag behöver den i morgon.
Jag behöver mer tid.
Jag behöver nycklarna.
Jag behöver skölja munnen.
Jag läser spanska.
Jag studerar spanska.
Jag vill städa huset innan mina föräldrar kommer tillbaka.
Framtiden tillhör inte de ängsliga, den tillhör de modiga.
Hon är vår granne.
Våren är här.
Våran har kommit.
Våren är kommen.
Det där var en utmärkt putt.
Jag har fått nog!
Jag bor här.
Vad lagar du?
Stanna!
Ingen vet.
Jag äter här.
Din hund är här.
Er hund är här.
Han är på väg att gå.
Den är väldigt stor.
Mig vantar kort.
Först till kvarn får först mala.
Jag älskar äpplen.
Ett stort tack för din hjälp.
Ett stort tack för er hjälp.
Grattis på födelsedagen!
Varför gjorde han det där?
Varför gjorde han så?
Vad heter den här gatan?
Kärleken är blind.
Jag ska lära dig hur man spelar schack.
Min dröm är att leva fredfullt i byn.
Jag brukade spela tennis.
Jag spelade tennis.
Många vackra blommor blommar på våren.
Enligt hans åsikt, ja.
Min pappa är inte hemma just nu.
Hon varnade barnen för att leka på gatan.
Det här är en vän till mig.
Jag skulle vilja ha en flaska hostmedicin.
Jag skulle vilja hyra en bil.
I fjol var april den varmaste månaden.
Jag heter Henry.
Herregud, jag kommer komma för sent till lektionen.
Ursäkta mig, talar du engelska?
Hon har ännu fler böcker.
Hon har solglasögon.
Hon gillar att springa.
Hungrig?
Jag litar på dig.
Jag litar på er.
Jag är hungrig eftersom jag inte åt frukost.
Det finns blott ett alternativ.
Grekiska är inget enkelt språk.
Grekiska är inget lätt språk.
Du är en idiot.
Håll käften!
Vissa studenter kommer inte att komma tillbaka nästa termin.
Några studenter kommer inte att komma tillbaka nästa termin.
Tack för er gästfrihet.
Tack för din gästfrihet.
Bron var byggd av romarna.
Bron byggdes av romarna.
Mannen vaknar.
Den rosa kudden är ren.
Den nuvarande regeringen har många problem.
Den korta kvinnan har på sig en svart kostym.
Strumporna luktar illa.
Läraren och eleverna är i museet.
Den unga mannen är läkare.
Det här landet heter Ryssland.
Detta är min lärare. Han heter herr Haddad.
Tvätta dina händer.
Välkommen hem till oss!
Välkomna hem till oss!
Vad tänker du på?
Vilken färg är din hår?
Vilken färg har ditt hår?
Vilken frukt är röd?
Vad har du i din påse?
Vad är växelkursen?
Mr. Smith kom.
Jag besöker honom varannan dag.
Du verkar ha förväxlat mig med min storebror.
John bryr sig inte ett dugg om sina kläder.
Så vitt jag vet är han inte lat.
Vi tittade alla ut genom fönstret.
Vi drack soju i karaokebaren.
Jag förstår mig inte på musik.
Kan du skicka saltet?
Spanska är hans modersmål.
Jag har stängt alla sex fönster.
Jag vet egentligen inte.
Jag vet inte riktigt.
Var är tvättrummet?
Han var modig.
Hur många minuter blir det om du omvandlar 48 timmar till minuter?
Ja.
Man kan lära sig många ord genom att läsa.
Solen är röd.
Det här är min fru, Edita.
Han stängde dörren.
Ingenting kan inte existera, för om det gjorde det så skulle det vara någonting.
Katten är på mattan.
Sockret är inne i påsen.
Jag blöder om knät.
Jag kan inte Svenska.
Jag pratar inte svenska.
Jag talar inte svenska.
Jag talar inte tyska.
Ingen bryr sig om vad du tycker.
Våren är här.
Ställ den var som helst.
Min mor nynnade för sig själv medan hon stökade på med matlagningen i köken.
Gillar du att äta fisk?
Jag måste bege mig nu.
Jag måste gå nu.
Jag måste bege mig nu.
Kan du se det där?
Skål!
Vilken lång gurka!
Vi behöver en ambulans.
Hatten är din.
Han älskar tåg.
Nej, inte riktigt.
Han borde avslöja alltihop och möta konsekvenserna.
Jag vet inte vad det är.
Varför behöver du de här pengarna?
Varför behöver du dessa pengar?
Jag är egentligen en universitetslärare.
Jag hittar inte det jag vill ha.
Det är läggdags.
Trevligt att träffas.
God dag.
Jag är kär i dig.
Det är risk att du blir en rejäl karl.
Räcker tiotusen yen?
Sluta att bita på naglarna.
Jag har ont i fötterna.
Det går fint!
Varför går inte människor i ide?
Han gräver sin egen grav.
Det är bara en dröm.
Jag kom hit i går.
Jag fick ett brev från min vän.
Vi har två barn.
Jag är arg.
Jag är för gammal för den här världen.
Jag gör det om de betalar mig.
Sluta upp med det omedelbart.
En vän i handen är bättre än tio i skogen!
Kan du inte ge me lite pengar?
Gnugga fläcken med vinäger.
Hon är inte ung längre. Hon är åtminstone 30 år gammal.
Men när jag försökte vrida duschkranen rann en svart, bubblig vätska ut.
Jag heter Farshad.
Att förstå dig är verkligen riktigt svårt.
Jag vill ha fem köttbullar.
Du har spillt lite ketchup på din slips.
Han låg på rygg.
Han har en bil.
Han bor inuti ett äpple.
Sådant är livet.
Är du Japansk?
Vad gjorde du med den här boken?
Vad gjorde du av den där boken?
Du borde inte vara arg.
Fråga mig någonting enklare.
Jag lyssnar på Björks senaste låt.
Får jag gå på toaletten?
Vart ska vi gå?
Du kan gå.
Du borde gå.
Den där dunkudden ser dyr ut.
Hon bestämde sig för att säga upp sig från sitt jobb.
"Den gamle och havet" är en roman av Hemingway.
Presidenten har avskaffat slaveriet.
Stäng din bok.
Stäng er bok.
Stäng igen din bok.
Stäng igen er bok.
Jag kan springa lika snabbt som Bill.
Jag är ledsen, jag tror inte att jag kommer kunna.
Jag åker dit varje år.
Vilken stor hund!
I går var det torsdag.
Mitt skosnöre fastnade i rulltrappan.
Hantverkaren lovade att komma nästa dag.
Allt gick bra.
Min mor sade åt mig att uppföra mig.
Jag talar japanska väl.
Tala högre så att alla kan höra dig.
Hur mår din mor?
Hur mår din mamma?
Glöm henne.
När man talar om trollen.
Det blir tre euro.
Himlen och helvetet existerar i mans hjärtor.
Vad är haken?
Kort hår passar henne verkligen.
Jag gillar verkligen inte Apple-produkter.
Jag oroar mig inte så mycket om mitt CV.
Ingen är för gammal för att lära sig.
Inga stjärnor syntes på himlen.
Har brevbäraren redan kommit?
Efter söndag kommer måndag.
Hon har en ödletatuering på låret.
De fångade räven med en fälla.
Var är chefen?
Den andra delen av boken utspelar sig i England.
Hon hjälpte dem med bagaget.
Det här är en turkisk tradition.
Det här är en väldigt tidsödande uppgift.
Jag är en vegetarian som äter massor av kött.
Jag har förlorat min PIN-kod!
Jag växte upp med att titta på Pokémon.
De övertalade mig att stanna ett tag till.
Wikipedia är den bästa encyklopedin på nätet.
Drick inte så mycket öl.
Vad kostar en öl?
Torka dina tårar.
De här är pojkar och de där är flickor.
Envar har rätt till skydd för de moraliska och materiella intressen, som härröra från varje vetenskapligt, litterärt eller konstnärligt verk, till vilket han är upphovsman.
Nästan tre.
Hunden är smart.
Jag har gått och tänkte på det hela dagen.
Jag har tänkt på det hela dagen.
Vissa fiskar kan ändra sitt kön.
Vissa fiskar kan byta kön.
Plastfolie är tillverkad i polyethylen.
En liten vinst är bättre än en stor förlust.
En liter mjölk innehåller ungefär trettio gram protein.
Frihet kostar.
Det fungerar inte.
Den fungerar inte.
Klava överförenklar allting.
Du kommer att få stå till svars för detta, Ibragim!
Var student har sin egen dator.
Varje student har sin egen dator.
Var elev har sin egen dator.
Varje elev har sin egen dator.
Vänta, skjut inte!
Is smälter i vatten.
Gjort är gjort.
Det var hans eget fel.
Vill du dansa med mig?
Jag heter Wang Jiaming.
Det här är mina byxor.
Jag behöver hjälp.
Översätt inte den här meningen!
Du tycker inte om mig.
Hur står det till? Jag har inte sett dig på evigheter!
Här är en mening, med stavelseantalet, som i en haiku.
Här är en mening, med stavelseantalet, som i en haiku.
Radion dog.
På tal om herr Tanaka, har du sett honom på sistone?
Jag är nöjd.
Jag är belåten.
Jag tycker inte om ägg.
Jag gillar inte ägg.
Jag ogillar ägg.
Han är en författare.
Det ska snöa idag.
Han studerar.
Han pluggar.
Vänta en stund.
Jag oroar mig över hans hälsa.
Han tappade kontrollen över bilen i kurvan.
Ät mer grönsaker.
De stal min vinflaska!
Storleken har ingen betydelse.
Varför hände det här?
Välkommen tillbaka. Vi har saknat dig!
Det erbjudandet låter för bra för att vara sant. Vad är haken?
Ditt hus är stort.
Ert hus är stort.
Han studerade hur fåglar flyger.
Jag har glömt min PIN-kod.
Det här svärdet är i gott skick.
Tror du på spöken?
Ta dig ett glas.
Ta en drink.
Vi är bekanta med den här sången.
Jag kommer aldrig att lämna dig.
Det finns ett parallellt universum i Bermudatriangeln.
Kommer du hit ofta?
Var är satelliterna?
Jag kunde svära på att någonting rörde sig.
Jag kände ett tryck på min axel och vände mig om.
Detta var en skön känsla.
Det här var en skön känsla.
Livet är orättvist.
Du förstör alltid allting.
En bild säger mer än tusen ord.
Jag kom hit tillsammans med mina vänner.
Det kommer att bli ganska kyligt.
De kommer från Sverige.
Du kommer från Sverige.
Kejsar Hadrianus lät bygga Hadrianus mur.
Han kan inte ha tappat bort sina nycklar.
Jag har köpt en bil.
Bomben exploderade för två dagar sedan.
Byggdes denna mur för att hålla människor ute eller för att hålla dem inne?
Byggdes denna mur för att hålla människor ute eller inne?
Byggdes den här muren för att hålla folk ute eller för att hålla dem inne?
Det rör mig inte i ryggen vad de säger.
Jag minns att jag mötte drottningen.
Hoppas medan du lever!
Det kommer inte göra ont.
Jag var på väg ut.
Men vad vill du?
Du har lättare för att komma ihåg saker än jag.
Jag hoppas att få se renar under min resa till Sverige.
Korrekt!
Det är sant.
Koka riset!
Den tillhör min bror.
Skämta inte med mig!
En kopp kaffe, tack.
Han gillar att springa.
Ge den till honom.
Ge det till honom.
Ge det till henne.
Ge den till henne.
Livet är ett uppvaknande efter ett annat.
En kopp kaffe, tack.
Jag kände mig lätt som en fjäder.
Peking är större än Rom.
Skulle du kunna förklara reglerna för mig, tack?
Skulle ni kunna förklara reglerna för mig, tack?
Ingendera är vacker.
Hon hittade jobb som maskinskriverska.
Skulle du vilja ha lite äggröra?
Talar du turkiska?
Det här är en rökfri kupé.
Behöver du hjälp med att bära något?
Behöver ni hjälp med att bära något?
Snabba er, ungar, annars missar ni skolbussen.
Zürich betraktas som en större finansiell knutpunkt.
Så du och Hanna planerar att gifta er?
Man bör läsa många böcker när man är ung.
Jag hatar dig väldigt mycket.
Var har hon lärt sig italienska?
Jag skulle vilja följa med, men jag är pank.
De skyndade sig till olycksplatsen.
Varför är himlen blå?
Jag bryr mig inte ett skit.
Jag kom på det.
Problemet är att pojken aldrig gör vad han blir tillsagd att göra.
Min bror har aldrig bestigit Mt Fuji.
Jag heter Jack.
Jag älskar min mamma.
Jag älskar min mamma.
Han är inte en av oss.
Han sade till henne att han älskade henne.
Flickan gick till skogen för att plocka svamp.
Kasta ingenting på marken.
Att ta genvägar sparar pengar på kort sikt men förlorar kunder på lång sikt.
Huvudstaden i Ukraina är Kiev.
Tre öl och en tequila tack!
Följer du med mig till affären?
Han är en gentleman.
Jag vill inte bo ensam.
Hon kommer kanske imorgon.
Huvudstaden i Ukraina är Kiev.
Jag tycker att vi ska vänta en halvtimme till.
Huvudstaden i Ukraina är Kiev.
Jag skulle vilja se dem igen.
Jag skulle vilja träffa dem igen.
Det finns många öar i Grekland.
Jag följer inte med.
Jag kommer inte på någonting.
Vad är det för fel på dig?
Hon kommer att betala för allting.
Min mor tycker mycket om té.
Vill ni ha té eller kaffe?
Jag bad honom att koka lite té.
Jag skulle inte vilja vara i hennes skor.
Han förblev obesegrad under hela sin karriär.
Hunden var upptagen med att gräva ner sitt ben i trädgården.
De flesta slott omges av en vallgrav.
Skratt smittar av sig.
Han sprang.
Han springer.
Det är min bok.
Hästen är min.
Jag skiter i vad du säger!
Jag har ingen kommentar.
Fem gånger sju är trettiofem.
Håll käften, annars åker du ut.
Folk som har varit med om så kallade 'lucida drömmar' beskriver dem ofta som 'verkligare än verkligheten'. De beskriver också verkligheten efter att de vaknat från en 'lucid dröm' som 'en nyckfull dröm'.
Han bor i Kyoto.
Hon bor i Kyoto.
Vad är skillnaden mellan en duva?
Seansdeltagare försöker få kontakt med de döda.
Hon befann sig på platsen för brottet.
Hon var på brottsplatsen.
Var är du nu?
Jag tycker om inte den här platsen.
Jag gillar inte den här platsen.
Jag tycker inte om det här stället.
Jag gillar inte det här stället.
Hur löser jag det här problemet?
Hur löser jag detta problem?
Tom är en duktig cricketspelare.
Är du rädd för skräckfilmer?
Är du rädd för rysare?
Det här är Carrie Underwoods senaste album.
Tom vill inte bli läkare, trots att han är väldigt på naturvetenskap.
Bränslenivån är under tom.
Tom samlade på kaffekoppar.
Föredrar du en manlig eller kvinnlig doktor?
Han går upp tidigt.
Han stiger upp tidigt.
Han kliver upp tidigt.
Jorden är där vi alla bor.
Tom hade tur som hittade sina nycklar.
De här skorna passar perfekt.
Det finns ett brev för dig.
Vi ska se en utländsk film ikväll.
Ungefär 9,4% av jordens yta är täckt av skog.
Hade du roligt i helgen?
Många människor litar inte på regeringen.
Jag hatar alla slags insekter.
Tom dömde en konsttävling.
Planet har nyss lyft.
Min katt hade ihjäl en ekorre.
Min mormors sjuksköterska är väldigt snäll.
Min farmors sjuksköterska är väldigt snäll.
Bajkalsjön i Ryssland är världens djupaste sjö.
Någon tappade sin plånbok.
Någon tappade en plånbok.
Marknaden öppnar klockan nio på morgonen.
Äter du kött eller är du vegetarian?
Äter ni kött eller är ni vegetarianer?
Jag protesterade när kyparen försökte ta min tallrik.
Vår värd erbjöd oss en drink.
Tom kan köra gaffeltruck.
En dag skulle jag vilja äga en segelbåt.
Hur många böcker äger du?
Tom hade ingen anledning att vara arg.
Mor stannade i bilen medan far handlade.
Mamma stannade i bilen medan pappa handlade.
Datorreparationen tog hela dagen.
Jordens måne är en naturlig satellit.
Våren är min favoritårstid.
Den ekonomiska situationen är inte bra just nu.
Väggarna i det gamla huset var inte raka.
Jag avskyr att se djur lida.
De gick mot porten.
Vi planerar en resa till New York.
Det är Marys tur att diska.
Varje morgon läser jag om vädret i tidningen.
Läraren välkomnade de nya studenterna.
Trottoarerna var blöta efter regnet.
Miljoner vilda djur lever i Alaska.
Många använder uttagsautomater för att ta ut pengar.
Tom undrar om det är sant.
Vädret är sämre i dag än i går.
Ett år senare föddes Paul.
Kor äter gräs.
Var köpte du denne klänning?
Var är ingången?
Vem sjunger den här sången?
Du har rätt. Jag tar en taxi.
Är det vad du vill?
Jag kommer inte ihåg vad hon heter.
Jag minns inte hennes namn.
Rökning dödar.
Om ett mänskligt liv är konvext, kan vi optimera det.
Kassören stoppade kundens varor i en påse.
Tack för ditt hårda arbete.
Tack för ert hårda arbete.
En förbipasserande bil körde i en vattenpöl och stänkte ned hela mig.
Jag behöver en kniv.
Behöver du pengar?
Behöver ni pengar?
Det är väldigt varmt idag.
Snart är det vår.
Han arbetar inte här längre.
Vi vet ingenting om honom.
Jag talar klingonska med dig.
Jag talar klingonska med er.
Jag föreslår honom till ordförande oavsett om du är för det eller inte.
Mödrar brukade säga till sina söner att om dom masturberade skulle dom bli blinda.
Russin är skrumpnade vindruvor.
Studerar eller jobbar du?
Jag äger två böcker.
Äh, tyst med dig.
Var är han?
Är det här franska?
Är det här franskt?
Är det här fransk?
Färglösa gröna idéer sover rasande.
Vi sätter julgranen här.
Vi ställer julgranen här.
Vad vill du köpa?
Koka lite vatten.
Jag orkar inte mer! Jag har inte sovit på tre dagar!
Jag arbetar 3 timmar varje söndagsmorgon.
Jag åkte till Italien för andra gången 1980.
Jag har att skynda!
Ut härifrån! Allihopa!
Glad mors dag!
Pappa är inte hemma.
Hunden är människans bästa vän.
Pojken var så trött att han inte kunde ta ett steg till.
Jag betalar med mitt kort.
Tvätta händerna innan du äter.
Har du tappat vettet?
Du är längre än mig.
När kommer du tillbaka?
Visa mig var Puerto Rico är på kartan.
Jag säger det till dig för sjuttioelfte gången – Nej!
Jane ger aldrig vika.
Jane prutar aldrig på sina anspråk.
Jane ger aldrig med sig.
Jag letar efter mina nycklar.
Någon satte dit honom.
Han är vid hennes sida.
Krig startar inte bara som vintern startar, utan snarare är det människor som startar ett krig.
Jag har inte tid för dig.
Jag har inte tid för er.
Vi vill att regeringen ska tjäna hela nationen.
Jag är vacker.
Jag är i bilen.
De äter inte kött.
De är vegetarianer.
Jag har inget emot att göra hushållssysslorna.
Jag tycker om att läsa innan jag går och lägger mig.
Du litar fullständigt på honom.
Ni litar fullständigt på honom.
Ubåten var tvungen att bryta igenom ett tunt istäcke för att kunna gå upp till ytan.
Vill du ha lite äggröra?
Kan du latin?
Finns det en tvättmaskin i huset?
Så romantiskt!
Det här är min häst.
Detta är min häst.
Jag älskar doften av papper när man slår upp en gammal bok.
Jag arbetar här.
Jag jobbar här.
Filosofi är egentligen hemlängtan; Längtan att vara hemma överallt.
Ett språk är en dialekt med en armé och en flotta.
Jag behöver ett frimärke.
Min kudde är så mjuk!
Jag är kvinna.
Jag känner inga blinda män.
Får jag också komma?
"Hur gammal är du?" "Jag är sexton år."
Han stiger upp klockan sju.
Jag missade tåget med bara några minuter.
Jag kan köra.
Jag har inte druckit kaffe än.
I morgon kommer jag inte att vara här.
Var så god och ge mig något att äta.
Hon drömde om vilda jaguarer.
Han är bara en amatör.
Han snarkade högt medan han sov.
Tre glassar, tack.
Han emigrerade till Australien.
En förbipasserande filmade polisens våld med sin mobiltelefon.
Människan uppfann atombomben, men ingen mus hade någonsin kommit på idén att konstruera en musfälla!
Mary har redan gått.
Jag tror hon är 40 år.
Vatten består av syre och väte.
Vad är klockan?
Han är min bror.
Jag lyssnar på musik.
Magsmärtorna är borta.
Kaniner gillar morötter.
Det är något med honom som jag inte gillar.
Det är någonting med honom som jag inte tycker om.
Skulle du kunna skriva ner länken till den sajten?
De gick tidigt.
Han kände sig trött.
Flygplanet ankommer klockan åtta.
Honom har hon inte sett på länge.
Hon har inte sett honom på länge.
Vi frågade honom vad han hette.
Jag har precis kommit tillbaka från Sverige.
Vi vill inte vänta längre.
Huset ligger vackert till.
Föraren körde om bilen.
Hon blev polis.
Jag tycker inte om honom, men jag gillar henne.
Hon har inte råd med det.
Han målar inte väggarna utan tapetserar dem.
Jag blev kär i dig.
Jag förälskade mig i dig.
Visade han dig bilden?
Den bilen är hans.
Varför ljuger du?
Varför ljuger ni?
Han kommer tillbaka sex.
Stillhet är guld.
Vad betyder "Tatoeba"?
Träffade du honom?
Jag gillar hundar och min syster gillar katter.
Jag tycker om hundar och min syster tycker om katter.
Pandor är väldigt smarta.
Varför är en del översättningar gråa?
Jag har skrivit ned alla siffror upp till trettioett.
Han kan inte utläsa vad det står på pappret.
De närmar sig.
Jar har ett hus i bergen.
Jag är rädd för bussen.
De har läst en intressant bok.
Det står bra till med min familj, tack.
Min familj mår bra, tack.
Jag går hem.
Jag har bröder.
Ja, så vitt jag vet.
Jag kan inte finna min flickväns klitoris.
Lyssnar du?
Det har varit ett dödsfall i din familj.
Detta är ett litet steg för en människa men ett jättekliv för mänskligheten.
Den tycker om att röka tobak.
Det tycker om att röka tobak.
Kan du inte skriva med kulspetspenna?
Jag kan inte.
En gång i tiden trodde man att människor inte kunde flyga.
Knivspetsen är vass.
Hon har stora bröst.
Jag skulle vilja åka till Frankrike någon gång.
Du kan skriva på vilket språk du vill. På Tatoeba är alla språk jämlika.
Jag tappade tålamodet.
"Du, min herre, är en imperialist!" "Och du, min herre, är ett troll!"
Jag studerar konsthistoria.
Mina vänner stod vid min sida under rättegången.
Mina vänner svek mig inte under rättegången.
Fler och fler studenter ansluter sig till protesterna.
Jag vill kunna läsa japanska.
Jag struntar hellre i skolan och spelar tv-spel istället.
Jag är ingen häxa.
Jag är orolig för honom.
Han bad om min hjälp.
Är du jänkare?
De vägrade låta tågen röra på sig.
Det dom sökte var en man som han själv.
De stödde honom och hans politik fortfarande.
Detta innebar att de var för svaga för att orsaka mer problem.
De krävde stränga straff för de södra rebellerna.
Han slutade aldrig att skriva.
Han dömde Brown till hängning.
Han besökte ett barnhem i Texas.
Han flydde från teatern efter mordet.
Han verkade trivas med sitt liv och sitt arbete.
Han hörde illa och kunde inte gå.
Finns du?
Finns vi?
President Truman var tvungen att fatta ett svårt beslut.
President Truman var tvungen att ta ett svårt beslut.
Importen av brittiska varor ökade.
Britterna trodde att amerikanerna överträdde deras lag.
Britterna tyckte att amerikanerna överträdde deras lag.
De allierade kontrollerade alla större irakiska städer.
Det var ett extremt grymt krig.
Många ryssar krävde ett slut på kriget.
Det är inte söndag varje dag.
Ingen gjorde något annat än att dansa.
Ingen vet säkert hur många människor som dog.
Alla pratade om det.
Republikanerna var rasande.
Jag vill inte ha era hus.
Jag vill inte ha dina hus.
Valet låg mycket nära.
Turkiet var starkare än Grekland.
Våldet varade i två veckor.
Nixon var på väg att bli president.
Al Smiths föräldrar kom från Irland.
Det rådde brist på importerad olja.
President Grant har inte gjort något olaglig.
1891 blev Liliuokalani Hawaiis drottning.
Kung George tog kontroll över kolonin 1752.
Han har glasögon.
Ormen frestade Eva.
Jag dödade Gud.
Jag har trott på Kylie Minogue sedan 12 juni 1998.
Jag mutade polisen.
Jag behöver kompisar.
Hur går det, sötnos?
Skriv under på den sprickade linjen.
Eftersom jag hade träffat honom en gång förut, kände jag igen honom direkt.
Eftersom jag hade träffat honom en gång innan, kände jag genast igen honom.
Låt oss hoppas att hon kommer.
Hörde du klickljudet?
Du är gammal nog att förstå.
Du är tillräckligt gammal för att förstå.
Vem talar?
Vem pratar?
Jag föddes sådan här!
Den här cd kostar tio dollar.
De gjorde en märklig upptäckt.
Jag visste att jag var tvungen att berätta sanningen för honom, men jag kunde inte förmå mig till det.
Jag kan inte göra det ogjort.
Terrorism är den viktigaste faktorn för delningen av ett land och skapandet av självständiga regioner.
Jag hatar dig.
Det var en så kraftfull explosion att taket flög av.
Får jag lov?
Det är säkert att äta fiskarna.
Det är säkert att äta fisken.
Om du inte studerar mer så kommer du helt säkert att misslyckas.
Vilka skolor härstammar från det Buddistiska tänkandet?
Dörrar är inte så dåliga som du tror.
Trots att jag har läst engelska 6 år i skolan talar jag det inte bra.
Mark stöter på allt som rör sig.
Den första gruppen studerar på morgonen, den andra på kvällen.
Det värsta med sommaren är värmen.
Det värsta med sommaren är hettan.
Ett bra vin behöver inte annonseras.
Hinner du?
Jag ser inget!
Jag har ingen katt.
Jag har beslutat mig för att svara på alla frågor offentligt.
Denna byggnad håller på att rasa samman.
Max förklarade för Julia varför han inte kunde komma på hennes avskedsfest.
Jag kan inte hjälpa dig.
Jag kan inte hjälpa er.
Jag talar lite skotsk galiska.
Hans förklaring var inte tillräcklig.
Det är det som är kruxet.
Smakar mjölken från den här renen verkligen gott?
Jag spelar ofta volleyboll.
Nästan alla hundar lever.
Vad kostar en öl?
Hej allihopa!
Jag är mycket trött.
Hon talar ryska.
Din fråga har inget svar.
Er fråga har inget svar.
Jag har svårt att tro på det.
Peking förändras så fort.
Det här är inte min åsikt, bara min översättning!
Jag använder Twitter.
Jag har lagat radion åt honom.
Förlåt för att jag stör, men min bil är trasig, skulle du kunna hjälpa mig?
Kossan säger "mu", tuppen säger "kuckeliku", grisen säger "nöff, nöff", ankan säger "kvack, kvack" och katten säger "mjau".
Du måste återbetala dina skulder.
Ni måste återbetala era skulder.
Många har samlats.
Pojken hoppar.
Hästen hoppar.
Flickan hoppar.
Hunden hoppar.
Vem läser?
Vem är det som läser?
Två barn sitter på staketet.
Du frågar fel person.
Min hund skäller hela tiden.
Det låter som en bra idé.
Gissa vem som kommer i kväll.
Att filosofera är att lära sig dö.
Är vädret fint?
Är hon trevlig?
Jag ser huset.
Ulster har minst förluster av alla boxare i ligan.
Jag måste ha drömt det.
En kungs dotter är en prinsessa.
Överlappning kan inträffa.
Varför är de här?
Det spelas inte mycket fotboll där.
Jag talar lite spanska.
Hon talar portugisiska.
Jag gillar inte kvinnor utan personalitet.
Varför gjorde han en sån sak?
Alla äpplen som faller till marken äts upp av grisarna.
Kartan hänger på väggen.
Hur stavas det?
"Tammi" med två m. Alltså T-A-M-M-I.
Han har inga vänner.
Jag har lånat en bil.
Låna aldrig en bil.
Jag har lånat ett bord.
Jag har lånat två böcker.
Talar du svenska?
Pratar du svenska?
Ja, lite grand.
Nej, inte alls.
Nej, jag förstår dig inte.
Tack, jag förstår nu.
Var finns det en telefon?
Finns det en busshållplats här i närheten?
Ja, där borta.
Kan du säga mig hur man går till amerikanska ambassaden?
Kan jag få köpa några vykort?
Jag skulle vilja köpa några vykort.
Hur många vill ni ha?
En krona och femtio öre.
Hur mycket blir det?
Det blir fyra kronor, tack.
Vi äter lunch.
Vi äter middag.
Vi äter frukost.
Kan jag få se på matsedeln?
Kan jag få se på menyn?
Kan jag få ett par ostsmörgåsar?
Skulle jag kunna få ett par ostsmörgåsar?
Vad vill ni ha att dricka? Kaffe?
Skulle jag kunna få ett glas mjölk, tack?
Kan jag få ett glas vatt?
Skulle jag kunna få ett glas öl, tack?
Skulle jag kunna få ett glas vin, tack?
Lite smör och bröd.
Det finns en restaurang här.
Det finns en buss här.
Det är en buss här.
Det finns en krona här.
Det är en krona här.
Det finns en telefon här.
Det finns en smörgås här.
Det är en smörgås här.
Det finns en hållplats här.
Det finns en busshållplats här.
Det finns ett vykort här.
Det står ett glas här.
Det finns ett glas här.
Det är ett par här.
Det finns ett par här.
Det finns ett hotell här.
Finns det en telefon här?
Jag talar svenska.
Jag pratar svenska.
Greta går till ambassaden.
Greta går till ambassaden.
Du ska tala svenska.
Du kommer att tala svenska.
Ni ska tala svenska.
Ni kommer att tala svenska.
Du ska tala svenska.
Du kan förstå svenska.
Ni kan förstå svenska.
En kopp kaffe kostar en krona.
Kostar en kopp kaffe en krona?
Herr Berg hjälper dig.
Hjälper du fröken Hansson?
Du vill hjälpa mig.
Jag hjälper dig.
Jag hjälper dig.
Jag ska hjälpa dig.
Jag ska hjälpa dig.
Jag kommer till hotellet.
Jag vill komma till hotellet.
Ett bi surrar.
Tittar de på oss?
Jag tror att jag äntligen ska pensionera mig.
När han åker till Europa kommer han att besöka många museer.
Ge mig en av dina bilder, tack.
Dr. Georges sekreterare är japanska.
Spinoza var en panteist.
Hör du mig bra nu?
Det finns mjölk i kylskåpet.
Jag önskar att jag vore ung igen.
Vem uppfanns telefonen av?
Det är hälsosamt att vara galen.
De gick och fiskade i går.
Hon föreslog för honom att resa utomlands medan han fortfarande är ung.
Hon rådde honom att ta medicinen.
Hon frågade honom varför han grät.
Hon slog ihjäl honom med en golfklubba.
Hon bet honom.
Hon lyckades inte övertala honom till att hålla tal.
Hon försökte inte att översätta brevet.
Hon lurade honom.
Hon gav honom en massa pengar.
Hon har känt honom länge.
Hon hatar honom.
Hon hörde honom sjunga.
Hon hjälpte honom.
Hon hjälper honom.
Hon slog honom.
Hon kramade honom.
Hon sparkade honom.
Hon kysste honom på pannan.
Hon kysste honom.
Hon vet bättre än att argumentera med honom.
Hon gillar honom.
Hon älskar honom.
Hon saknar honom.
Hon beordrade honom att städa upp sitt rum.
Hon övertalade honom att göra det fastän hon visste att det inte var en god idé.
Hon kvävde honom med en kudde.
Hon såg fram emot att gå på bio med honom.
Hon väckte honom.
Ingå i en överenskommelse med mig och bli en ung magisk flicka!
Telefonen är trasig.
Jag talar spanska med Gud, italienska med kvinnor, franska med män och tyska med min häst.
Sen sjöng jag en dum låt om en myra som försökte brottas med ett tuggummi.
Jag köpte en grön soffa igår, men den gick inte in genom dörren, så jag fick lämna tillbaka den.
Det där måste vara historiens rödaste finne.
Jag såg på när de flådde en människa den dagen.
Han är min bror, inte min far.
Jag vill dö med Getter Jaani.
Och slutligen, tolv poäng till Estland!
Är din mor hemma?
Han kan inte ens skriva sitt eget namn.
Det finns mer än 4000 språk i världen.
Det finns mer än 4000 språk i världen.
Hur dags gick du och lade dig igår?
Kan jag använda telefonen?
Jag har stånd.
Man gör leksaker i den här fabriken.
Jag gillar verkligen hårdkokta ägg.
Hur ofta äter du fisk?
Jag är på ett gräsligt humör i dag för jag har inte tillräckligt med pengar.
Vladivostok är en stad i Ryssland.
Och varför frågar du?
Vad oroar du dig för?
Medan han pratade hördes ljudet av ett skott som avlossades.
Medan han pratade hördes ett skott avlossas.
Vår galax heter Vintergatan.
Grattis på födelsedagen.
Det är bara en tidsfråga.
Många träd tappar sina löv på vintern.
Många träd tappar löven på vintern.
Till min förvåning var han bra på att sjunga.
Det finns ett akut behov av bloddonationer.
Jag tror det är dags för mig att dra.
Skynda dig tillbaka.
Spring!
Vilken är din favoritsvordom?
Vilken nagellack är din favorit?
Vilket är ditt favoritnagellack?
Vilken är din favoritprotestsång?
Vilken är din favoritsuperhjälte?
Vem är din favoritsuperhjälte?
Det regnar idag. Var är mitt paraply?
Det här är inte min åsikt, bara min översättning!
Han ljuger.
Vad säger han?
Det var oförlåtligt.
Det är vad alla säger.
Du älskar kaffe.
Vi har diskuterat det här problemet nyligen.
Magdalena och Ania är goda vänner.
Både Magdalena och Ania är från Polen.
Nuförtiden verkar alla vara lyckliga.
Stanna gärna kvar efter konserten. Vi kommer signera autografer.
Tímea är en ungrare som bor i Polen.
Medtävlanden tjuvstartade två gånger.
Han behöver en stege.
Jag har varit död förr, och det var inte så illa.
Den största skillnaden mellan bandy och innebandy är att bandy spelas på is.
Koreaner tycker inte om koriander.
Varför alltid jag?
Min pappa är starkare än din.
När jag väl öppnade ögonen igen satt Amina och stirrade på mig genom botten av sitt ölglas.
Vad heter den här gatan?
Grodan och jag turades om att gissa vad det hemliga receptet var.
Jag köpte inte den där boken.
Vem är din lärare?
Min vän George ska till Japan i sommar.
Vet du vem hon är?
Mitt hus ligger i norra delen av staden.
Snälla, förlåt mig.
Kvinnan är naken.
Många unga romare åkte till Grekland.
Låt oss berätta allt vi vet.
Två gånger sju är fjorton.
Att mingla med folk på fester kan vara förskräckande för blyga människor.
Jag hittade ett väldigt trevligt ställe i går.
Läs inte denna mening.
Tråkar jag ut dig?
Mår du bra?
Tycker du att jag är ful?
Tycker ni att jag är ful?
Gråt inte.
Har du ätit?
Har du någonsin varit på TV?
Hur är det med din pappa?
Hur mår din pappa?
Hur länge måste jag stanna här?
Hur många självmord tror du att det sker varje år i Japan?
Hur var din dag?
Hur var din kväll?
Jag åt för mycket.
Jag sa inte att det inte var okej att äta.
Jag avskyr att ha med kräsna barn att göra.
Jag kunde inte föreställa mig att jag skulle känna såhär för dig.
Jag försökte att inte gråta.
Jag undrade bara om du har lyckats hitta någonstans att bo.
Jag försöker bara tjäna en slant.
Att äta en klyfta vitlök varje dag, är det nyttigt för dig?
Är det bra för hälsan att äta en vitlöksklyfta om dagen?
Är det nyttigt för dig att äta fisk?
Är det moraliskt fel att äta kött?
Min hund åt min läxa.
Var snäll och stäng av motorn.
Det fanns mycket som vi helt enkelt inte hade tid att göra.
Det står en man med en pistol i handen i dörren.
Det står en man med en pistol i handen vid dörren.
Den här ordboken kan komma till användning.
Vi älskar dig så mycket.
Vad krävs för att man ska få lite hjälp?
Vad gör du idag?
Din engelska är grammatiskt riktig, men ibland låter det du säger bara inte som något en modersmålstalare skulle säga.
Din engelska är grammatikalisk, men ibland låter det som du säger bara inte som någonting som en modersmålstalare skulle säga.
Han sa att han inte visste.
Han sa att han inte vet.
Inget är omöjligt för Gud.
Mannen är naken.
Vi älskar picknickar.
Inatt var det väldigt varmt och kvavt och jag sov inget vidare.
På två drag kommer Kasparov att ställa motståndaren i schack.
Du måste förbereda dig för det värsta!
Hon är orolig över din säkerhet.
Hon är orolig över er säkerhet.
Det var i det huset som jag föddes i.
Han är en hjälte.
Sådan är lagen.
Vi är lika inför lagen.
Tror du att Steve Jobs skulle ha varit lika framgångsrik som han varit om hans efternamn varit "Joobs" istället?
Jag vet inte när han kommer, men när han gör det, kommer han att göra sitt bästa.
Jag kan inte gå förrän han kommer.
Och så förälskade sig lejonet i tackan.
Är du okej?
Du borde inte döma folk efter utseendet.
Man ska inte döma folk efter utseendet.
Detta är en häst.
Den här hunden är min.
Det är kvavt här inne.
Det är kvalmigt här inne.
Kan du släppa av mig vid biblioteket?
Kom in och sitt ner, är du snäll.
Att lära sig koreanska är svårt.
Varför köpte du en blomma?
Russin är torkade vindruvor.
Jag reser ofta.
Det är regn på väg.
Det är ingen leksak!
Du måste sluta ljuga för dig själv.
Han blir lätt trött.
Jag läser den här boken.
Egentligen inte.
Båda gick till fönstret för att titta ut.
Jag måste sova.
Han är konstig ibland.
Jag öppnade asken. Den var tom.
Vad är det för fel på mig?
Jag är finsk.
Han är ett matematiskt geni.
Jag är jättetjock.
Tom tog bussen till skolan.
Tom tog ut en penna och började skriva.
Tom tog fram en penna och började skriva.
Tom tog av sig rocken eftersom det var för varmt för att ha den på sig.
Tom tog av sig rocken och kastade den på golvet.
Tom tog av sig sin rock och sina handskar.
Tom tog av sig sina kläder och gick in i duschen.
Tom verkar sova.
Tom sa att han ville komma bort från stan ett tag.
Tom sade att han ville komma bort från staden ett tag.
Tom räddade hunden ifrån att bli uppäten av de hungriga soldaterna.
Tom slutade röka.
Tom behöver köpa en ny regnrock.
Tom gjorde många misstag.
Tom ser väldigt glad ut.
Tom lever ur hand i mun.
Tom är inte den gitarrist som han brukade vara.
Tom är inte lång.
Tom är inte här.
Tom är inte en bra kock.
Tom är den perfekta fadern.
Tom är verkligen ledsen.
Tom kommer aldrig i tid.
Tom är vänsterhänt, men han skriver med höger hand.
Tom kommer också till festen.
Tom kan komma på vår fest i morgon.
Tom är en mycket stark man.
Tom är en hemmaman.
Tom har två söner. Båda av dem bor i Boston.
Tom har två sönder. Bägge bor i Boston.
Tom har för mycket arbete att göra.
Tom har tre onklar.
Tom har något i sin hand.
Tom har haft problem med sitt vänstra öga sen olyckan.
Tom har studerat franska i ungefär tre år.
Tom har redan druckit tre koppar kaffe.
Tom tar en promenad varje eftermiddag.
Tom samlade ihop alla sina saker.
Tom gjorde klart läxan innan kvällsmaten.
Tom somnade till slut.
Tom äter som en gris.
Tom arbetar inte lika hårt som han brukade.
Tom vet inte vart han skall gå.
Tom vet inte vad han ska beställa.
Tom kommer inte överens med sina grannar.
Tom känner inte för att prata just nu.
Tom dricker inte.
Tom tycker inte om huset han bor i.
Tom försvann utan att lämna ett spår.
Tom försvann utan ett spår.
Tom visste inte vad han skulle göra härnäst.
Tom visste inte vad det var meningen att han skulle göra.
Tom gjorde det för skojs skull.
Tom bestämde sig för att säga upp sig.
Tom kunde inte bestämma sig.
Tom kunde inte bestämma sig omedelbart.
Tom kunde inte hitta någon att prata med.
Tom kunde inte besvara en endaste fråga på gårdagens test.
Tom kollade datumet.
Tom kan inte läsa utan glasögon.
Tom kan inte bestämma sig för vilken kamera han ska köpa.
Tom kom för att be oss om hjälp.
Tom kom hit för att be oss om hjälp.
Tom kom hit för att be om vår hjälp.
Tom ringer mig nästan varje dag.
Tom åt en handfull russin.
Tom bär alltid en karta och kompass i sin väska.
Detta är min vän Tom.
Allt är Toms fel.
Jag tvivlar på att Tom är glad.
Jag tvivlar på att Tom är lycklig.
Tom undrade om det som Mary sade var sant.
Tom brukade hata Mary. Nu älskar han henne.
Tom tackade Mary för hennes råd.
Tom skrattade sällan åt Marys skämt.
Tom låtsades inte förstå vad Mary sa.
Tom missade chansen att åka till Boston med Mary.
Tom fick Mary att gråta.
Tom skrattade åt Mary.
Tom skrattade åt alla Marys skämt.
Tom vet Marys hunds namn.
Tom kysste Mary på pannan.
Tom dödade Mary.
Tom kan bara inte komma överens med Mary.
Tom är granne till Mary.
Tom är trogen Mary.
Tom är Mary trogen.
Tom är förlovad med Marys lillasyster.
Tom förlät Mary på hennes dödsbädd.
Tom känner inte att han kan lita på Mary.
Tom tvivlar inte på Marys förmåga att utföra jobbet.
Tom kunde knappt förstå vad Mary sade.
Tom ser Mary som en hjältinna.
Tom tror att Mary fattade rätt beslut.
Tom blev trött på att alltid behöva betala notan varenda gång han gick ut med Mary.
Tom bad Maria att öppna fönstret.
Tom bad Mary hålla ett tal.
Tom frågade Mary om hon kunde hjälpa honom.
Tom och Mary vaknade tidigt för att se årets första soluppgång.
Tom och Mary paddlade kanot längs med floden sist jag såg dem.
Tom och Mary verkar inte hungriga.
Tom och Mary verkar inte vara hungriga.
Tom och Mary avskyr varandra.
Tom berättade för Mary om John.
Om du vill vara fri, försttör då nu din TV.
Han har en vit katt.
Får jag öppna en burk?
Hur kan jag lösa det här problemet?
Hur kan jag lösa detta problem?
Tatoebaprojektet, som återfinns online på tatoeba.org, går ut på att skapa en stor databas med exempelmeningar översatta till många språk.
Jag ber om ursäkt för det sena svaret.
Vem är jag? Var kommer jag från? Finns det liv efter döden? Vad är meningen med livet på jorden?
Olyckligtvis släppte Tom ut katten ur säcken.
Det förklarar varför dörren är öppen.
Det förklarar varför dörren står öppen.
Hon läser tidningen varje morgon.
Du behöver inte vänta till slutet.
Klockan var nästan 2:30 när Tom till slut kom hem.
Det här är mannen som jag letat efter.
Jag är ingen nazist.
Kan du skicka mig den där grunkamojen?
Jag ville inte spendera mer tid på att arbeta med det där projektet.
Storebror ser dig.
Tom har en liten paj.
Jag antar att vi borde gå nu.
I begynnelsen skapade Gud himmel och jord.
I begynnelsen skapade Gud himmel och jord.
En katt är inte en person.
Jag ställer alarmklockan så att jag inte kommer för sent till jobbet imorgon.
Min bror är lärare.
Varför gör du så mot mig?
Hunden blöder.
Det här är första gången jag skriver ett brev på spanska.
Ingen rök utan eld.
Nordkoreas tillbakadragne ledare besöker Ryssland för förhandlingar om energi.
Jag tror att jag är utarbetad.
Jag tror att jag är överansträngd.
Jag vet inte vad rätt svar är.
Kan du inte röra dig fortfarande?
Bladen är gula.
Var är äpplen?
Amy, du borde gifta dig med honom.
Mina väskor är packade.
Han beskrev i detalj vad som hade hänt.
För tillfället har jag inte nog med pengar.
Tyskland ligger mitt i Europa.
Det finns regler att följa.
Den här filmen är för barn.
Skriv endast ut jämna sidor, tack.
Kan du tala kinesiska?
Kan du prata kinesiska?
Kan du kinesiska?
Jag tycker inte om dig längre.
Vi litar på honom.
Har du pojk- eller flickvän? Var träffade du hen?
Har du pojk- eller flickvän? Var träffade du honom eller henne?
Helga är ett svenskt namn.
Jag ville bli astrofysiker en gång i tiden.
Hur länge kommer det här kalla vädret att hålla på?
När såg du senast Tom?
Vad har du för bevis på att det var Tom som stal din mors halsband?
Toms nya skjorta krympte i tvätten så nu passar den inte.
Toms bil är lätt igenkännbar eftersom det är en stor buckla i den främre stötfångaren.
Tom undrade varför Mary var så sen.
Tom var tokförälskad i Mary.
Tom vill att Mary ska träffa hans mor.
Tom ville hämnas.
Tom försökte sälja sin gamla videobandspelare istället för att slänga den, men ingen köpte den, så det slutade med att han slängde den.
Tom trodde att ingen var hemma.
Tom verkar inte vilja sänka priset.
Tom säger att han aldrig har försökt äta hundmat.
Tom sa att han trodde att Mary fortfarande bodde hos sina föräldrar.
Tom låtsades inte veta vart han skulle gå.
Tom lämnade tv:n på hela natten.
Tom har dörrarna låsta om natten.
Tom vet verkligen inte vad han ska göra.
Tom är van att ta snabba beslut.
Tom är ute.
Tom är en främling i den här staden.
Tom har inget lokalsinne.
Tom har aldrig sett Mary så arg.
Tom gick vilse.
Tom satte sig i förarsätet och körde iväg.
Tom kände sig väldigt ensam.
Tom tror inte att detta är någon tillfällighet.
Tom gillar inte Marys attityd.
Tom tycker inte om Marys attityd.
Tom ville inte berätta för Mary att han hade förlorat alla hennes pengar.
Tom tänkte inte på det.
Tom förväntade sig inte riktigt att Mary skulle svara på hans fråga.
Tom gav inte upp.
Tom fick inte något gjort idag.
Tom visste inte var han skulle börja.
Tom borde definitivt ha fått dödsstraff.
Tom bestämde sig för att skjuta upp beslutet.
Tom kunde inte kontrollera sig själv.
Tom kunde knappt gå.
Tom är verkligen snål.
Tom behöver sannerligen inte mer pengar.
Tom verkar inte komma åt sina data.
Tom verkar inte komma åt sin data.
Tom kan inte bestämma sig för vad han ska köpa.
Tom kan skriva med båda händerna.
Tom kan tala flytande franska.
Tom kan tala franska flytande.
Tom kan prata flytande franska.
Tom kan prata franska flytande.
Tom bad om en filt och en kudde.
Tom och Mary har varit gifta i tre år.
Tom klagar nästan aldrig på någonting.
Jag hade aldrig kunnat gissa att Tom och Mary skulle bli kära i varandra.
Jag tror att det är osannolikt att Tom kommer till festen själv.
Hur länge har du känt Tom?
Hur länge har ni känt Tom?
Du behöver koppla av.
Någon förstörde min kamera.
Någon gjorde sönder min kamera.
Någon hade sönder min kamera.
Jag vill inte prata om det.
Jag sa att jag var förvirrad.
Jag är korean.
Jag äter ett äpple.
Tom tycker inte om den här färgen.
Pojkarna och flickorna leker i trädgården.
Gud skapade jorden på sex dagar.
Den här pojken är lat.
Jag har ett par med päron.
Hoppa!
När jag springer, blir jag svettig.
Jag ska till Paris.
Hur såg rånaren ut?
Han är trött på mina problem.
Förlåt.
Jag är från Brasilien.
Svarta katter betyder otur.
Slåss som en man!
Vi ses i morgon!
Min far var ett träd.
Kontakta henne om du har några frågor.
De betedde sig underligt.
Du missbrukar dina maktbefogenheter.
Vi har en begränsad budget.
Jag är höjdrädd.
Vi hade rätt.
Vad är det för fel på honom?
Hon har vackra ögon.
Hon är kvart över nio.
Talaren är ung.
Det verkar som att Taro inte har några tjejkompisar.
Hon är inte vackrare än deras mor.
Min dator har hängt sig.
Han höll på att bli en känd sångare.
Hon är stark.
Jag kokar fortfarande råriset.
Jag är inte för trött.
Jag väckte dig.
Jag tycker inte om det.
Jag tycker inte om det där.
Jag gillar det inte.
Jag gillar frukt.
Jag tycker om frukt.
Behöver du dricka vin?
Behöver ni dricka vin?
Du är vårt enda hopp.
Är han från Japan?
Är hon Japansk?
Ge mig dina tankar.
Skitsamma.
Jag har fått nog.
Låter det bekant?
Mina föräldrar är väldigt stränga.
Det kan jag inte utesluta.
Jag med.
Du är trygg här med mig.
För att dölja det faktum att hon var en princessa förklädde hon sig till en pojke och flydde från slottet.
Jag vill inte gifta mig.
Jag har aldrig träffat dig i verkligheten.
Det var inget sammanträffande.
Nunnorna sjunger.
Det är en harpa.
Jag blödde näsblod idag.
Det är Babas röst.
Det är en gammal kvinnas röst.
Min syster tycker om Ultraman.
Papegojan är död.
Dags att sticka.
Vad kämpar du för?
Han är en drama queen.
Mjölk är en vanlig dryck.
Jag går till arbetet varje dag.
Jag promenerar till jobbet varje dag.
Tro på dig själv.
Var snäll mot andra.
Din önskan har gått i uppfyllelse.
Är det din egen idé?
På inrådan av sina astronomer bestämde sig Alexander den store för att inte attackera Egypten och for till Indien istället.
Jag är i San Diego och ni bara måste komma och hälsa på mig!
Utsikten är fantastisk.
Du borde komma och hälsa på oss!
Ni borde komma och hälsa på oss!
Det är roligt att spela baseball.
Alkohol löser inga problem, men det gör inte mjölk heller.
Han gråter alltid när han är full.
Han säger att han älskar blommorna.
Jag kan bo i gästrummet.
Det finns nästan inget syre i rummet.
Det var ett oförlåtligt misstag.
Jag åt med min lillebror.
Bron förbinder de två städerna.
Igår eftermiddag skrev jag ett brev.
Du måste ha blandat ihop mig med någon annan.
Min fru slår mig.
Matade du papegojorna?
Minns du den gången vi åkte till Paris?
Vi hade en överenskommelse. Du bröt den.
Har du lite bröd? Jag ska mata duvorna.
Jag tycker om att mata duvorna.
Hon äter inte kött, eller hur?
Vi kysstes.
Det är en papegoja i fågelburen.
Män vet inget om kvinnor.
Vi har ett väldigt allvarligt problem.
Jag är fortfarande arg på henne.
Det trodde jag aldrig om dig.
Det är första min far skrev.
Gör vad du vill.
Du har bara en chans att svara rätt.
Han hade snö upp till knäna.
Jag är finsk, men jag talar svenska också.
Jag vill inte laga mat.
Jag har inte tid att laga mat.
Vilken är din favoritsnabbmatsrestaurang?
Vilken är din favoritsnabbmatsrestaurang?
Vilken är din favoritsnabbmatsrestaurang?
Vilken är din favoritsnabbmatsrestaurang?
Jag har aldrig varit i Argentina.
Snabbmat kan vara beroendeframkallande.
Har du pengarna?
Du är anhållen.
Jag gillar utmaningar.
Det finns inga droger här.
Ett land utan horhus är inget land.
Se dig omkring.
Är det etiskt att ge honom intervjufrågorna i förväg?
Välkommen till mitt liv.
En diskret hyllning till olycksoffren hölls igår.
Skaffa dig ett liv.
Må balroger äta dig.
Du är fin i håret.
Var hälsad, gillesbroder.
Bara kärlek kan krossa ditt hjärta.
Bara kärlek kan krossa hjärtat.
Bara kärlek kan krossa ens hjärta.
Endast kärlek kan krossa ditt hjärta.
Endast kärlek kan krossa hjärtat.
Endast kärlek kan krossa ens hjärta.
Han låtsas vara döv.
Vilken är nästa station?
Kommer han hem klockan sex?
Hur var det?
Flickan dricker te.
Han talar lite engelska.
Jag äter med händerna.
Han hade ont i huvudet.
Hur kan jag få dig att ändra dig?
Det här börjar bli svårt.
François, är denna din?
François, är detta ditt?
Hur länge tänker du stanna här?
Han tycker mycket om musik.
Det är länge sedan jag såg honom.
Vem gick du med?
Jag blev avskedad.
Tom var klädd helt i svart.
Tom var helt hjälplös.
Tom stängde av tv:n.
Tom tycker att det är tillräckligt bra.
Det är bäst att du inte väntar längre.
I det mest spännande ögonblicket, såg alla väldigt spända ut.
Hur är det möjligt?
Hos dig eller hos mig?
Hon är envis.
Allt var väldigt bra.
Droppe blod.
Det är ett rökmoln över landskapet.
Det är ett rökmoln över provinsen.
Det här företaget är listat på Parisbörsen.
Tom dyker oftast upp i tid.
Tom såg Mary på TV.
Tom lurade dig.
Tom fick slut på bensin.
Tom skalade potatis.
Så du ska ingenstans imorgon?
Det är ett gammalt manuskript.
Jag kan inte engelska.
Du har inget bra minne.
Jag hatar politik.
Jag kan springa.
Hon är ungefär i min ålder.
Hon älskar katter.
Jag är säker.
Hon blandar ofta ihop socker och salt.
Nu du kommer till Frankrike ska vi åka till Marseille.
Gårdagen är historia. Morgondagen är ett mysterium. Dagen idag är en gåva. Det är därför den kallas för nuet.
Förlåt honom om du kan. Han är oskyldig.
Jag beordrade ungarna att vara tysta, men de fortstatte att väsnas.
England och Skottland är grannar.
Jag har bara sett det en gång.
Jag har bara sett den en gång.
Snart är det din tur, Bashar!
Marias hår är långt.
Håll utkik efter en skallig och svettig kille.
Du måste vara Tim Norton.
Hur kan ni inte gilla honom?
Hur kan ni inte tycka om honom?
Hur kan du inte gilla honom?
Hur kan du inte tycka om honom?
Jag är ingen läkare.
Hon gråter alltid när han är full.
I min värld är alla en ponny, som äter regnbågar och bajsar fjärilar.
Jag är ingen läkare.
Många vet inte om att antibiotika är verkningslösa mot virussjukdomar.
Varför är du så trött?
Du behöver bara be om det.
Ni behöver bara be om det.
Ni behöver bara be om den.
Du behöver bara be om den.
Ingenting spelar egentligen någon roll.
Jag uppskattar verkligen din hjälp.
Det påminde mig om dig.
Det påminde mig om er.
Jag vill sova lite längre.
Du hade läst.
Katten satt på mattan.
Jag är inte din slav.
Vet du hur hans far dog?
Mamma, var är toalettpappersrullen?
Kinesisk filosofi är bäst.
Hon är grym.
Jag fattar.
Jag har bott sex månader i Kina.
Jag skulle vilja ha ett svar.
Du borde verkligen sluta röka.
Fastän det låter märkligt är det sant det hon sade.
Han sover under dagarna och jobbar under nätterna.
Många fiskar dog.
När PC-fel saktar ner dig, vad kan du göra ?
Plutonium-239 har en halveringstid på 24 100 år.
43-åriga kvinna misstänks ha skjutit ihjäl sin make.
Naturen är full av mysterium.
Städerskan trodde att hon bara gjorde sitt jobb - i själva verket förstörde hon ett modernt konstverk värt miljoner. Nu brottas museet med hur det ska hantera krisen.
Det här spelet är baserat på en roman.
Det är din rättighet.
Ut ur mitt hus!
Vi ses vid huset!
Under soffan finns många dammråttor.
Det finns många dammråttor under soffan.
Du är guld värd.
Jag får åksjuka.
Det var en bra dag.
Barn dricker mer vatten, äter mer mat och andas mer luft per kilogram kroppsvikt än vuxna.
Efter avslutat samtal sä­­ger han vänligt adjö och önskar mig en trevlig kväll.
De kommer att ha jättekul.
Han fick jobbet.
Jane slutade samla på nallar vid tjugo års ålder.
Där tar du troligen fel.
Var är dina nycklar?
Jag drog mig ur.
Det är en film som alla borde se.
Min mamma lagar mat åt mig.
Döda havet lever. Det lockar turister från världens alla hörn.
Skulle ni kunna ta en titt på mitt första inlägg och berätta vad ni tycker om det?
Behovet av reformer i Italien är enormt.
Vilken årstid gillar du mest, våren eller hösten?
De är inte alltid där.
Det är en oklar historia.
Jag har glömt mina glasögon.
Var har du gömt julklappen?
Var det inte Kafka som skrev att en bok måste bli yxan för det frusna havet inom oss?
Jag såg du-vet-vem i dag på torget.
Krokodilarna har vassa tänder.
Krokodiler har vassa tänder.
Middagen var toppen.
De älskar varandra väldigt mycket.
Jag gillar den personen.
Jag förlorade allt.
Han går fort.
Hon dukade av bordet efter middagen.
Jag känner mig lättare än luft.
När jag öppnade dörren hade jag sönder låset.
Det här är mitt rum.
Det fanns lite dagg imorse.
Min mormor bodde hos oss.
Hon är upptagen.
Vi måste skjuta upp vår avresa.
Jag tror inte det blir bättre än så!
Du måste läsa mellan raderna.
Man måste läsa mellan raderna.
Det gör inte så ont.
Gammal är äldst.
Gör honom inte besviken.
Vill någon ha en öl?
Upp med händerna! Detta är ett rån.
Du kan gå om du vill.
Ni kan gå om ni vill.
Hotellet har en hemtrevlig atmosfär.
Följ den bilen.
Jag var hemma.
Låt mig betala.
Jag var tvungen att ge upp.
Jag fick ge upp.
Jag fick säga upp mig.
Jag var tvungen att säga upp mig.
Tatoeba var tillfälligt otillgängligt.
Han är på sjukhuset.
Hon är online flera timmar varje dag.
"Kebabmorden" verkar ha lösts.
Han är inte sjuk.
Tack för alla dina kommentarer!
En bok är tunn och den andra är tjock; den tjocka har cirka 200 sidor.
Du luktar så gott.
Han gick långsamt så att barnet kunde följa med.
Han gick långsamt så att barnet kunde hänga med.
Han gick långsamt så att barnet kunde hinna med.
Han gick sakta så att barnet kunde hinna med.
Han gick sakta så att barnet kunde hänga med.
Han gick sakta så att barnet kunde följa med.
Han gick långsamt så att barnen skulle kunna klara av att följa efter.
Han har ett stort hus och två bilar.
Han studerade hårt så han inte skulle misslyckas.
Han litar mycket på sin assistent.
Han verkade besviken över resultaten.
Han säger alltid elaka saker om sin fru.
Han är väldigt smart, så alla gillar honom.
Han tänkte att det skulle vara vettigt att acceptera erbjudandet.
Han behövde inte ta med sig ett paraply.
Det var inte nödvändigt att han skulle ta med ett paraply.
Ofta kommer han inte till skolan.
Han visade mig hennes bild i smyg.
Han visade mig hennes foto i smyg.
Han visade mig hennes fotografi i smyg.
Han har ingen chans att återhämta sig.
Det finns ingen chans att han kommer att återhämta sig.
Han gick ut ur rummet så fort som jag gick in.
Han kan inte ha sagt något så dumt.
Han gillar musik mycket.
Han älskar musik.
Han gillar verkligen musik mycket.
Han lät mig sova över en natt.
Han var sjuk, så han kunde inte komma.
Han är vänligt mot alla sina klasskamrater.
Han spelade golf varje dag under semestern.
Han gick in på banken utklädd som en vakt.
Han gick ut ur rummet utan att säga ett ord.
Han försökte att göra sin fru lycklig, men han kunde inte.
Han gick vilse när han var ute och gick i skogen.
Han övar på att spela gitarr tills sent på kvällen.
Han vann första pris på schackturneringen.
Han har vanan att läsa tidningar under måltider.
Hur lärde du dig att spela fiol?
Jag kommer känna mig ensam när du har gått.
Hur länge kommer det här kalla vädret att fortsätta?
Hur hände trafikolyckan?
Det han sa visade sig vara en lögn.
Oavsätt hur mycket hon äter, så går hon aldrig upp i vikt.
När jag kom hem, upptäckte jag att jag hade tappat bort min plånbok.
John fick Mary att hoppa till.
John fick Mary att hoppa.
Jag dricker alltid två koppar kaffe varje morgon.
Premiärministern kommer att hålla en presskonferens imorgon.
Jag tror att jag skall köpa en ny bil.
Jag är inte säker på när han kommer att komma.
Jag har hört den låten sjungen på franska.
Jag har hört den franska versionen av den här låten.
Jag ville ringa några telefonsamtal.
Jag kommer förklara incidenten.
Låt mig berätta för dig om fallet.
Jag kommer att vara sexton år gammal på min nästa födelsedag.
Jag tycker att hon är en ärlig kvinna.
Jag tyckte att den här filmen var väldigt intressant.
Jag lånade ut en del pengar till min vän.
Jag gjorde ett dåligt misstag på provet.
Jag gjorde ett allvarligt misstag på provet.
Jag begick ett allvarligt misstag på provet.
Jag tycker att du behöver tänka på framtiden.
Jag tycker att du borde tänka på framtiden.
Jag var inte medveten om att du mådde så dåligt.
Jag var inte medveten om att du mådde så dåligt.
Jag tycker att han är en skicklig person.
Jag tycker att han är skicklig.
Jag vet inte hur man spelar golf överhuvudtaget.
Jag kunde inte gå på hans födelsedagskalas.
Jag höll i repet hårt så att jag inte skulle falla.
Jag höll hårt i repet så att jag inte skulle falla.
Jag är säker på att jag kommer vinna tennismatchen.
Jag kände mig väldigt lättad när jag hörde nyheterna.
Jag översatte dikten så gott som jag kunde.
Jag tycker att det är tragiskt att inte ha några vänner.
Geologen klev in i limon.
Lyssna!
Ja, sa hon, du har rätt.
Är jag fadern?
Hon är min fru.
Försöker du stöta på mig?
Hon är van vid att sitta.
Hur kommer det sig att du alltid är sen?
Hon skadades i en bilolycka.
Herre, var nådig mot min son, ty han är epileptiker och lider fruktansvärt därav, för han faller ofta in i elden, och ofta ner i vattnet.
Rökning kan orsaka impotens.
Hon sjunger otroligt bra.
Fyratusen meningar kan översättas på ett år av en talande man.
Jag måste gå på min kusins dop.
Känner du igen honom?
Den som är född i Sverige är svensk.
Jag känner mig så vacker.
Grönt står för hopp.
Paris är en ganska dyr stad.
Jag lär mig språket själv.
Det kommer inte att fungera.
Det kommer inte att funka.
Det kommer inte att gå.
Han är så söt.
Jag har en känsla av att hon kommer att komma idag.
Jag ska arbeta under sportlovet.
Jag ska plugga engelska i eftermiddag.
Jag ska studera engelska i eftermiddag.
Jag ska ta med min son till djurparken i eftermiddag.
Jag ser fram emot sommarlovet.
Jag börjar tappa tålamodet.
Jag vet inte om han är en doktor.
Jag vet inte om han är en läkare.
Jag kan inte hitta Tom. Har han redan gått?
Skala äpplet innan du äter det.
Hitta katten.
Hon dog av törst under torkan.
Det stör mig att hon alltid är sen.
Jag vill dansa.
Jag läser.
EU grundas för att få slut på de blodiga krigen mellan grannländerna, som gång på gång hade orsakat så mycket mänskligt lidande och till slut ledde till andra världskriget.
Jane låtsades alltid att hon var väldigt rik.
Från och med 1950 börjar en rad europeiska länder samarbeta ekonomiskt och politiskt för att bevara freden.
1950-talet karakteriseras av ett kalla krig mellan östblocket och västmakterna.
Det gjorde mig ytterst glad.
Hon rådde honom att prata om sitt liv i Förenta Staterna.
Frihetsgudinnan är symbolen för USA.
Vi träffades en vinter.
Jag är emot det.
Vi har sett henne.
Var ligger Mississippi?
Han drack öl.
Han drack en öl.
Vi spelar schack. Jag har redan tagit fyra av hans pjäser.
Använder du aftershave?
Använder ni aftershave?
Vissa kvinnor rakar inte benen.
Vissa kvinnor rakar inte sina ben.
Somliga kvinnor rakar inte benen.
Somliga kvinnor rakar inte sina ben.
Vad skulle ha veta?
Hon blev tvungen att förlita sig på sin inre styrka.
Jag vill samma svärdet som det!
Hon log åt mig medan hon sjöng en sång.
Ibland förstår jag mig inte på honom.
Ibland förstår jag inte honom.
Ibland förstår jag honom inte.
Vilken sport tycker du mest om?
Här är jag född och uppvuxen.
Bussen är tom, och ändå sätter han sig bredvid mig.
Franskan utvecklades från latin.
Jag har precis ätit färdig.
Vi har en reservation klockan halv sju.
Jag har levt här under en lång tid.
Jag känner mig väldigt förrådd.
Han är DJ.
Vad betyder katakres?
Stäng dörren! Det drar.
Soldaterna är döda.
Jag kom hem sent.
Tom och Mary hade kuddkrig.
Toms föräldrar bor i en gammal husvagn.
Staden var öde.
Vad heter hon nu igen?
Jag har en massa arbete att göra imorgon.
Han kommer alltid att älska henne.
Han återvände hem efter att ha varit borta under tio månader.
Vargar brukar inte attackera människor.
Jag behöver gå ner i vikt, så jag håller på med en diet.
Hon hjälpte den gamla mannen över vägen.
Han visade mig en massa vackra bilder.
Han visade mig massor av vackra bilder.
Jag kan inte komma ihåg den låtens melodi.
Den gamla kvinnan gick upp för trappan med möda.
När man har fått in en dålig vana, så är det inte enkelt att bli av med den.
Jag är på åttonde våningen.
Jag ska inte göra illa dig.
Årets icke-ord 2011 är "Kebabmord".
Håll bollen med båda händerna.
Jag är rädd för hundar.
Jag är nyfiken.
Rätta mig om jag har fel.
Det verkar som att jag har en lätt förkylning.
Förlåt att jag har orsakat dig så mycket besvär.
Hon håller på med en diet.
Hon är frånvarande för att hon är sjuk.
Han är tre år äldre än hon.
Han är tre år äldre än henne.
Hon vill veta vem det var som skickade blommorna.
Hon är nyfiken på att få reda på vem det var som skickade blommorna.
Jag vet inte exakt när jag kommer att komma tillbaka.
Jag skjuter upp min resa till Skottland tills det blir varmare.
Klockan är redan elva.
Hon kommer förmodligen.
Jag är överraskad att du vann priset.
Det är svårt att förstå hans teori.
Det är upp till dig att bestämma om vi skall gå eller inte.
Jag sa till henne en gång för alla att jag inte skulle gå och handla med henne.
Om inte den där gitarren vore så dyr, så skulle jag kunna köpa den.
Jag vill ha en båt som kan ta mig långt härifrån.
Det kommer försätta dig i fara.
Kaniner har långa öron och korta svansar.
Han har bott på det där hotellet de fem senaste dagarna.
Hon har inte varit i skolan på fem dagar.
De är på god fot med sina grannar.
Vi har gått runt hela sjön.
Du borde ha avvisat ett sådant orättvist förslag.
Det där är varför han blev arg.
Det där är anledningen varför han blev arg.
Stranden är ett idealiskt ställe för att barn att leka.
Det ligger en bok om dans på skrivbordet.
Vilka språk talas i Amerika?
Vilket land är störst, Japan eller England?
Hon hade precis börjat läsa boken när någon knackade på dörren.
Vart i Turkiet bor du?
Du jobbar för hårt. Ta det lugnt en stund.
Du går inte upp lika tidigt som din syster, eller hur?
Du ser precis ut som din storebror.
Du borde inte säga såna saker när barn är i närheten.
De senaste medicinska framgångarna är anmärkningsvärda.
Han la boken på hyllan.
Han tjänar tre gånger så mycket som jag.
Han tjänar tre gånger så mycket som jag gör.
Han tjänar tre gånger så mycket som jag.
Han tjänar tre gånger så mycket pengar som jag gör.
Han tjänar tre gånger så mycket pengar som jag.
Han berättade sin livshistoria för mig.
Tiderna förändras, och vi förändras med dem.
Mary försökte trösta Tom.
Att oroa sig är som en gungstol; det ger en någonting att göra men leder ingenstans.
Burj Khalifa är världens nuvarande högsta skyskrapa.
Vilken tid passar dig?
Vilken tid passar er?
Mary gillar att festa.
Det verkar som att Mary är full igen.
Tom är en desertör.
Tom är en värnpliktsvägrare.
Mary kände sig utstött.
Tom ville inte göra något han skulle komma att ångra.
Filmen inspirerades av boken med samma titel.
Jag sov som en stock.
Vad pratar hon om?
Depression är vanligt bland unga vuxna som har Asperger syndrom.
Mary är konstig.
Finns de?
Vi håller kontakt.
Jag vill inte prata om henne.
Varför bestämde du dig för att prata om det nu?
Jag tror inte att hon skulle förstå det.
Jag antar att han kommer tillbaka snart.
Rapporten ansågs vara falsk.
Vill ni att jag skall koka kaffe?
Min far fick mig att tvätta bilen.
Cowboy hoppade snabbt ut genom fönstret.
Ölglaset är nästan större än dig.
Kossan muar, tuppen galer, grisen grymtar, ankan kvackar och katten jamar.
Tom är plastikkirurg.
Jag är van vid att äta ensam.
Jag känner mig gammal.
Det påstås att det snart kommer ett val.
Den mannen dog av lungcancer för en vecka sedan.
Den kvinnan har två väskor.
John har en bil från Japan.
Jag gav tiggaren alla pengar jag hade.
I morgon är det jul.
Soldaten slog samman klackarna.
Den nya telefonboken är här!
Alice sover i mitt rum.
Du måste lyckas där dom största hjältarna har misslyckats.
Det var hans tystnad som gjorde henne arg.
Han vann allt.
Om du vill, så ring mig på eftermiddagen.
Hon heter Irina.
Jag trivs verkligen i Georgia.
Jag trivs verkligen i Georgien.
Hon gillade poesi och musik.
Jag önskar dig lycka.
Jag önskar dig allt väl.
Jag önskar dig lycka till.
Hon är fortfarande minderårig.
Jag läste att Brasiliens president är en kvinna. Hon kallas Dilma.
Jag läste att Brasiliens president är en kvinna. Hon kallas Dilma.
Du är lat!
Ni är lata!
Man stöter på japanska turister överallt.
Han har inte lyckats än.
Jag behöver köpa frimärken.
Jag glömde att ringa Herr Ford.
Du borde slå upp det ordet.
Du borde slå upp det ordet.
Vad tror du hände här?
Vad tror ni hände här?
Korsningen där olyckan inträffade ligger här i närheten.
Målet var offside.
Var är ingången?
Hade jag vetat skulle jag ha sagt det till dig.
Hans far vigde sitt liv åt vetenskapen.
Det är en skugga.
Jag kan inte stoppa blödningen.
Du sa att du var lycklig.
Ni sa att ni var lyckliga.
Deras favoritämne var eskatologi.
Jag lyssnar nästan aldrig på radio.
"Han har varit sjuk." "Jaså, jag hoppas att det inte är någonting allvarligt."
Han är någonstans i parken.
Sann kärlek existerar inte.
Jag kommer börja gråta!
Jag kommer börja grina!
Det har gått tre år sedan vi gifte oss.
Torka byxorna på elementet.
Jag hatar när mina kläder luktar cigarettrök.
Tom klarar sig jättebra.
Tom klarar sig mycket bra.
Jag köpte många böcker.
Jag köpte en massa böcker.
Vilken blomma som helst går bra, så länge den är röd.
Tom har bevisat att det fungerar.
Tom har bevisat att den fungerar.
Tom har bevisat att det går.
Herr Wang kom till Japan för att studera japanska.
De fulla sjömännen har ställt till med elände inne i baren.
Tom är en naturlig atlet.
Han låtsas.
Idag är det imorgon vi oroliga igår.
Tom är ett äckel.
Hon kom inte innan två.
Doktorn sa till herr Smith att sluta röka.
Mary är ganska orolig.
Mary är ganska stökig.
Var tålmodig.
Ha tålamod.
Var tålmodiga.
Tom kommer inte att göra det.
Hon sa själv att hon inte skulle bli kär i någon igen.
Han satt i stolen.
Han hjälper inte till hemma.
Jag sitter och studerar på biblioteket.
Det är din först arbetsuppgift.
Han är på tåget.
Alice har fantastiska benen.
Tom är en korgosse.
Tom är sångare i gosskör.
Varför följer du efter mig?
Varför förföljer du mig?
Varför förföljer ni mig?
Varför följer ni efter mig?
Det är 48 sjömän på skeppet.
Det är fyrtioåtta sjömän på skeppet.
Tom är neurolog.
Tom är nervspecialist.
Är det där franska?
Om du får någon tid över, använd den och gör dina läxor.
Tom är en kommunist.
Tom är en präst.
Sluta anmärka på Tom.
Sluta hacka på Tom.
Hur är ditt liv som gift?
Hur är ert liv som gifta?
Varför är tåget sent?
Varför frågar du mig?
Hur kom du dit?
Hur tog du dig dit?
Hur ska du klara dig?
Hur ska ni klara er?
Klä på dig fort.
Klä på er fort.
Vilken station är det här?
Vilken station är detta?
Hur klarar du det?
Hur lyckas du?
Jag behöver en cigarett.
Ska vi fika?
Det är inte en bra idé.
Jag tar en promenad.
Jag skulle vilja förbättra min franska, men Jag får inte tid med.
Vattenverket ligger inte långt från mitt hem.
Tom är en hippie.
Tom är en hipster.
Tom är en beatnik.
Vill du ha lite öl?
Jag har varit där mycket.
Alla studenterna i klassen gillar herr Smith.
Alla elever i klassen tycker om herr Smith.
Han kanske inte är ung.
Är du buddist?
Är du buddhist?
Det är hans julklapp.
Han satt alldeles tyst och tittade rakt fram.
De körde igenom flera samhällen på vägen.
Hon tittade på alla hus som gled förbi.
Hon undrar hur det se ut där de skulle bo.
Men allra mest undrade hon vad hette henne.
Då är jag framme.
Nå vad tycker di om mig?
Han lastade ur bilen.
Hon stängde försiktigt ytterdörren.
Så bullrig det var därinne.
Rummet verkar väldigt mörkt och kusligt.
Det ekade ödsligt.
De gick uppför trappan.
Jag letade efter mitt rum.
Du ska hitta dina leksaker och böcker.
Jag kände mig genast lite bättre.
Dessa fenomen inträffar, men sällan.
Vad är det för filtillägg?
England åker ut på straffar igen.
Aldrig prata med främlingar.
Vad gör tvättbjörnen i köket?
Hennes dröm är över.
Tom undrade vad Mary's efternamn kunde vara.
Transformation är födelse och död på en och samma gång.
Tom har inget perspektiv.
Vi värdesätter våra kunder.
Han skulle ha gjort det allaredan.
Han skulle ha gjort det redan.
Hon skulle ha gjort det redan.
Hon skulle ha gjort det allaredan.
Tom är sociopat.
Tom är oärlig.
Tom är bedräglig.
Tom är en flykting.
Tom är en rymling.
Tom är en landsflykting.
Tom är på väg.
Tom ryckte på axlarna.
De lät mig välja en present.
Tom studsade tillbaka.
Tom gjorde en bra putt.
Tom är en sportig typ.
Tom är en idrottare.
Tom är en idrottskille.
Esperanto talas i 120 länder runt om i världen.
Tom är kompetent.
Tom är skicklig.
Mary knäböjer.
Tom är en sympatisk kille.
Tom har dålig hygien.
Tom är blyg och feg.
Sätt i ett mynt.
Jag såg henne igår.
Jag såg henne i går.
Tom gick ut och dansade.
Tom är Marys skyddsling.
Tom är Marys protegé.
Tom såg förbryllad ut.
Tom såg villrådig ut.
Tom såg häpen ut.
Tom såg frågande ut.
Tom sjukanmälde sig.
Det var mitt nöje.
Tom blev avvisad.
Tom fick avslag.
Tom fick nej.
Tom fick korgen.
Tom är lång och smal.
Tom fritog gisslan.
Hennes hud var varm.
Titanic krockade i ett isberg.
Tom flämtade.
Tom flåsade.
Tom stönade.
Tom såg sig inte om.
Tom såg inte tillbaka.
Tom tänkte inte tillbaka.
Tom drog sig inte ur.
Tom backade inte ut.
Den här maten är glutenfri.
Tom säger att han är villig att göra det gratis.
Jag tror att jag kommer att kunna träffa dig snart.
"Är du svensk?" "Nej, schweizisk."
Hon gillade det.
Hon gillade den.
Hon tyckte om det.
Hon tyckte om den.
Tom är otrogen.
Tom är trolös.
Den är gjord av läder.
Den är gjord av skinn.
Åt du frukost?
Åt ni frukost?
Tom drack i tystnad.
Tom såg honom aldrig igen.
Det är gammal skåpmat.
Alice är min mamma.
Tom är en helbrägdagörare.
Vi blir inte yngre.
Vi blir inte yngre än så här.
Han är lagkapten.
Livet är inte lätt.
Japaner utbyter gåvor för att uttrycka sina känslor.
Tom bad mig om hjälp.
Något kommer att hända. Jag känner det på mig.
Visa oss runt.
Peka ut den.
Peka ut det.
Flytta på dig.
Det slutade bra.
Jag försöker komma på varför någon skulle göra något sådant.
Jag försöker komma på varför någon skulle göra någonting sådant.
Jag försöker komma på varför någon skulle få för sig att göra något sådant.
Jag försöker komma på varför någon skulle få för sig att göra någonting sådant.
Är det några frågor?
Vi ska inte på semester.
Det är ovanligt.
Jag fick dig.
Jag har dig.
Har du några syskon?
Tillsätt naturell yoghurt och sojamjölk.
Vi har problem.
Vi är i trubbel.
Vi är illa ute.
Vi är i knipa.
Vi har råkat illa ut.
Tom bestämde sig för att läsa juridik.
Jag tvättade bilen.
Jag ser fram emot det.
Det är för kallt.
Den är för kall.
Han är en väldigt hälsosam person.
Tror du att vi kommer att hitta hennes hus?
Tror ni att vi kommer att hitta hennes hus?
Detta är Ken. Han älskar sin hund.
Det här är Ken. Han älskar sin hund.
Vem sjunger den här sången?
När han kom hem, sov barnen redan.
Kvinnor känner att män ofta är väldigt komplicerade.
Om du inte vill dit, så åker vi inte dit.
Tom gjorde ett halv-färdigt jobb.
Det var en gång en kung som hade tre döttrar.
Nej, jag är engelsk.
Jag brukade simma i havet när jag var ett barn.
Nej, jag är engelsk.
"Är du svensk?" "Nej, jag är schweizisk."
Han har två bilar.
Bucklan var min.
Pottan var min.
Krukan var min.
Burken var min.
Kannan var min.
Grytan var min.
Haschet var mitt.
Det är min häst.
Jag är ledsen att jag har inte skrivit till dig på så länge.
Han har två bilar.
Tom kräver uppmärksamhet.
Tom har behov av uppmärksamhet.
Tom är en eldslukare.
Tuppen galer "Kuckeliku!" om morgonen.
Tack för senast.
Jag har skrivit ett brev.
Stormen sänkte temperaturen.
Han dog innan ambulansen kom.
Jag vill inte ha någon frukt.
Får den här lådan plats i skåpbilen?
Tom hade helt rätt.
Hon vill arbeta på ett sjukhus.
Såg du gårdagens avsnitt?
Jag föddes med tolv fingrar.
Jag gillar ris mer än bröd.
Hur länge ännu, Catilina, skall du missbruka vårt tålamod?
Hörde du det där?
Skolan är tråkig.
Det låter bekant.
Mary är en gold-digger.
När kom Susana tillbaka?
Köpte du läkemedlet?
De kallar den här planeten "Jord".
Du då, litar du på den här mannen?
Ni då, litar ni på den här mannen?
Jag ville träffa dig.
Jag vet att jag kommer att dö.
Du vet den där känslan?
De är svåra att hitta.
Anpassning är nyckeln till överlevnad.
Smaklökar är väldigt användbara.
Skynda dig!
Spring för livet!
Tom gillar reality-tv.
Tom tycker om reality-tv.
Du är inte rolig.
Du fattar inte, eller hur?
Ni fattar inte, eller hur?
En katt har en svans och fyra ben.
Måndag börjar på söndag.
Jag vill inte dö!
Jag har lucida drömmar.
Jag har klarsynta drömmar.
Jag har klardrömmar.
Det var bara en liten kärleksaffär.
Hon har små bröst, men jag har inget emot det.
Han sparkade honom medan han låg ner.
Tom bor med Mary i Memphis.
Hur tar jag mig till busshållplatsen?
Det är en encellig organism.
Jag har alltid varit en ensamvarg.
Det vet du inte.
Jag vill inte leva.
Tom lär sig engelska.
Tom stör Mary.
Tom håller på att somna.
Tom häller upp ett glas mjölk.
Tom masserar sina knän.
Tom masserar hans knän.
Spara lite glass åt mig.
Han är mycket förstående.
Men det är inte det sista tåget, eller?
Vi bakar kakor.
Skjut inte!
Varför vill du att världen ska känna till japanska trädgårdar?
Jag blandar majonnäs med ketchup.
Tuppen pickar på mitt ben.
Om du verkligen vill lyckas måste du tycka om att äta gift.
Våra gudar är döda.
Vet du var mina gamla glasögon är?
Det var poängen.
Mannen satte eld på sig själv.
Ser man på!
Ingen vill dit.
Jag behöver kaffe.
Kapitulera eller dö!
Hon bad sin lärare om råd.
Finns det någon som kan svara?
Är det någon som kan svara?
Säg någonting även om du inte vet rätt svar.
Vi kommer överens.
Vi kommer väl överens.
Du blir tvungen att laga mer mat.
Jag dödade en gud.
Jag bodde i det här huset som barn.
Ha ett bra liv.
Ha ett trevligt liv.
Ha ett bra liv.
Detta är första gången jag ber i en moské.
"Det är första gången jag river min ägare", sa katten.
De utgör att skickligt lag.
Vem brukade göra detta?
Vem brukade göra det här?
Det finns bara två primtal mellan 10 och 14.
Det är första gången jag parkerar min bil i skogen.
Det här företaget använder billig arbetskraft för att öka sina vinstmarginaler.
Jag är allergisk mot gluten.
Jag gör det för att jag måste.
Jag sade aldrig att det inte vad en bra idé.
Jag sa aldrig att det inte var en bra idé.
Ett enormt monster är på väg ned från berget.
Mary är nu en glad liten flicka.
Jag tog ut kakan ur ugnen.
Gör som jag!
Husen brinner.
Glöm inte att det finns undantag.
Vi tar kreditkort.
Om han inte går i skolan tänker jag inte prata med honom längre.
Tack för att du tröstade mig när jag var ledsen.
Förlusten av hennes far var väldigt smärtsamt för henne.
Kan du inte skriva "Pfirsichbäumchen"? Det är så simpelt.
Det är ett extremfall.
Jag har ingen aning om vad jag ska förvänta mig.
Jag skulle göra vad som helst för kärlek.
Jag skulle göra vad som helst för kärleken.
Stick!
Jag gillar inte huset.
Jag tycker inte om huset.
Jag gör det här för hennes skull.
Sluta vara så nyfiken.
Han blir rädd lätt.
Han blir lätt rädd.
Jag kan inte bullra. Barnet sover.
Min mamma jobbar på fabrik.
Hon går sällan, om någonsin, ensam på bio.
Jag ska till Paris i helgen.
Allting har ett pris, det goda visar sig vara dyrare än det onda.
Har du någonsin tvättat din bil?
Har ni någonsin tvättat er bil?
Ring brandkåren!
Vem håller du på?
Vem hejar du på?
Vilka håller du på?
Vilka hejar du på?
Har du grävt upp potatisar?
Är perfektion tråkigt?
Min syster har gett mig en iPhone, men jag vet inte hur man använder den.
Det startade en kedjereaktion.
Rör er inte!
Kan Tatoeba bidra till att rädda utrotningshotade språk?
Jag är inte din fru längre. Din fru är Tatoeba!
Var god, kryssa i den lämpliga rutan.
Det var en stor en.
"Vill du lämna ett meddelande?" "Nej, tack."
Visst är det möjligt om man vill.
Luften är fuktig.
Vänta!
Jag måste låna lite pengar.
Dayxa är min hustrus syster.
Dayxa är min svägerska.
Mohand är min halvbror.
Oroa dig inte. Han förstår inte tyska.
Oroa dig inte. Han kan inte tyska.
Den mänskliga handen har fem fingrar med naglar.
Det här är mitt skepp.
Vill ni spela tennis med oss?
Vill du spela tennis med oss?
Får jag raka av dina polisonger?
När kommenterade du en mening senast?
Han har inte på sig en hatt.
Han har inte på sig hatt.
Han har inte hatt på sig.
Han har inte en hatt på sig.
Han vet hur man flyger en helikopter.
Jag säger er, jag säger er, den Drakfödde kommer!
Det betyder slutet för ondskan, och för alla fiender av Skyrim.
Ty mörkret har passerat, och legenden gror ännu.
Är du ledsen?
Var ligger den svenska ambassaden?
Var finns det en svensk ambassad i USA?
Det finns en svensk ambassad i Washington D.C.
Var ligger den kinesiska ambassaden?
Var ligger den australiska ambassaden?
Var ligger den kanadensiska ambassaden?
Var ligger den danska ambassaden?
Var ligger den egyptiska ambassaden?
Var ligger den finska ambassaden?
Var ligger den grekiska ambassaden?
Var är den grekiska ambassaden?
Var ligger den ungerska ambassaden?
Var ligger den indiska ambassaden?
Var ligger den israeliska ambassaden?
Var ligger den italienska ambassaden?
Var ligger den nyzeeländska ambassaden?
Var ligger den norska ambassaden?
Var ligger den portugisiska ambassaden?
Var ligger den ryska ambassaden?
Var ligger den spanska ambassaden?
Var ligger den nederländska ambassaden?
Var ligger den turkiska ambassaden?
Var ligger den brittiska ambassaden?
Var ligger den amerikanska ambassaden?
Marys meningar är lätta att översätta.
Jag har korrigerat misstaget.
Ingen visste att du var i Tyskland.
Det är inte tillåtet för kvinnor att köra bil i Saudiarabien.
När kan vi mötas igen?
När kan vi träffas igen?
När kan vi ses igen?
Solen är vit.
Han är bög.
Jag vill leva i staden.
Nej, det här pappret är inte vitt.
Laurie älskar mig.
Nej, jag tittar inte på CNN.
Det är 99,9 procent effektivt.
Det är nittionio komma nio procent effektivt.
Vad är lufttemperaturen idag?
Han drack direkt från flaskan.
Han drack direkt ur flaskan.
Tom talade till Mary från den andra sidan.
Succé! Detta är den femtusende klingonska meningen på Tatoeba!
Många tror att fladdermöss är fåglar..
Många människor tror att fladdermöss är fåglar.
Det var hans beslut.
Jag älskar Lauries hår.
Han festar för mycket.
Vad vill du bli när du blir stor?
Varför skär du upp frukterna?
Hon måste vara död.
Han är rädd för katter.
De låter besvikna.
Du låter besviken.
Ni låter besvikna.
Hon har inga barn.
Ingenting är så enkelt som det verkar.
Inget är så enkelt som det verkar.
Jag tror du är svartsjuk.
Han är din vän.
Han är din kompis.
Hur använder man ätpinnar?
Jag ska presentera dig för några vänner som läser tyska.
Sophies finger blödde så mycket att blodet droppade ner på marken.
Jag skrev min första mening på tyska.
Jag skriver en mening på tyska.
Jag kan inte se dig.
Jag vet inte varför.
Jag vet inte vad jag vill.
Jag vill lära mig tyska med mina vänner.
Hon talar inte engelska.
Jag kommer att skriva en mening på tyska.
Jag ska skriva en mening på tyska.
Hans fru är svensk.
Det är min son.
Jag skriver korta meningar på svenska.
Jag skriver en sång på tyska.
Jag skriver en sång på tyska.
Jag skriver ett brev till min fru.
Jag räknar på tyska.
Jag läser det här brevet.
Algeriet ligger i Nordafrika.
Algeriet är mitt land.
Pfirsichbaeumchen är från Tyskland.
Jag lär mig svenska och tyska.
Du lär dig arabiska.
Var ligger Algeriet?
Jag ska precis till att skriva en mening på tyska.
Jag vill ha en bok på svenska.
Wenjin är en kinesisk kvinna.
En mans ansikte är hans självbiografi. En kvinnas ansikte är hennes skönlitterära verk.
Du såg hunden som tillhör den man som jag flirtade med.
Edward Sapir var en amerikansk lingvist.
Andorra är ett litet furstendöme beläget mellan Spanien och Frankrike.
Vad har hon gjort?
Mår han bra?
En man som kan två språk är värd två män.
Jag älskar Kalifornien.
Ingen är rik i mitt land.
Vi behöver dig.
Jag skriver en roman.
Vad skrev du igår?
Vill du ha någonting att äta?
Vill du ha något att äta?
Vill du ha nåt att äta?
Och om han har fel?
Hon är orolig för sin vikt.
Hon oroar sig för sin vikt.
Var snäll och påminn mig om jag glömmer bort.
Hennes syster bor i Skottland.
Det är precis som jag förväntade mig.
Hon är nästan sextio år gammal.
Ge mig ett halvt kilo äpplen.
De vill inte att du ska veta.
En tredjedel är mindre än en halva.
Var han fallskärmsjägare?
Varför bryr hon sig inte om mig längre?
Sverige heter "Sverige" på svenska.
Jag vill förändra världen.
Somalia heter "as-Sumal" på arabiska.
Syrien heter "Suriyah" på Arabiska.
Sverige är det största landet i Skandinavien.
En ponny är en liten häst.
Han ger ut böcker i Italien.
Den svarta kattungen hoppade för att undvika pölen, och passerade under den angränsande häcken.
Hur många århundraden finns det på ett millennium?
Hur många dagar gammal var jag när den här bilden togs?
Bor dem i Algeriet?
Han var riktigt kall.
Vad dom säger är sant.
Din cykel är mycket nyare än min.
Vi hinner inte i tid till mötet.
Dom bär dyrbara ringar.
De bär dyrbara ringar.
De bär dyra ringar.
Jag var väldigt glad.
Jag var mycket glad.
Vi översatte rapporten från engelska till afrikaans.
Jag kan faktiskt inte svaret.
Jag vet faktiskt inte svaret.
Tom åt någonting.
Tom har aldrig ätit rått hästkött.
Tom borde inte ha ätit så mycket.
Jag äter bara koscher mat.
Hur kom Tom in?
Hur tog sig Tom in?
Hur tog Tom sig in?
Tom låtsades inte höra Mary ropa hans namn.
Jag har ett tajt schema den här helgen.
Gå och byt om.
Frågade du Tom?
Tack så mycket.
Vad sa du till Tom?
Vad sa ni till Tom?
Vad berättade du för Tom?
Vad berättade ni för Tom?
Vad tycker du, Tom?
Jag kommer inte ihåg vilka artiklar jag har översatt och inte.
Jag översätter inte romaner längre.
Ta det lugnt.
Ta det i din egen takt.
Jag är inte din fiende.
Jag är inte er fiende.
Tom ser skräckslagen ut.
Varför är ni alla här?
Mary är där inne.
Jag fattar fortfarande inte.
Låt oss sköta vårt jobb.
Gör dig av med pistolen.
Få Tom att ringa mig.
Berätta för mig vad Tom sa.
Tom åt en snabb lunch.
Tom åt en snabblunch.
Tom åt en tidig middag.
Tom åt sig mätt.
Tom åt så mycket han orkade.
Tom åt upp ditt godis.
Tom äter ofta äggröra till frukost.
Jag kan inte bestämma var vi ska äta lunch...
Vänta en sekund.
Håll ett öga på Tom.
Hon är en ängel.
En man som inte spenderar tid med sin familj kan inte vara en riktig man.
Ge Tom allting.
Låt mig hämta Tom.
Låt mig prata med Tom.
Låt mig tala med Tom.
Håll dig borta från Tom.
Hälsa till Tom.
Ge mig din tröja.
Den tjocka tjejen äter för mycket sötsaker med mycket socker i.
Den tjocka flickan äter för mycket sötsaker med mycket socker i.
Det är väldigt intressant.
Han är flytande på Engelska.
Det fick mig att skratta.
Det är svårt att säga.
Hon var ung och oskyldig.
Oroa dig inte. Det är enkelt.
Oroa dig inte. Det är lätt.
Ödsla inte din tid.
Ödsla inte er tid.
Slösa inte bort er tid.
Slösa inte bort din tid.
Maska inte.
Slösa inte bort Toms tid.
Slösa inte Toms tid.
Rör inte dem.
Rör inte mina grejor.
Rör inte mina grejer.
Rör inte mina prylar.
Rör inte mina saker.
Tacka mig inte än.
Berätta inte för någon.
Prata inte med mig.
Tala inte med mig.
Ta inga risker.
Var inte uppkäftig.
Var inte kaxig.
Svara inte på det.
Få mig inte att döda dig.
Få mig inte att döda er.
Få mig inte att skada dig.
Tvinga mig inte att göra detta.
Tvinga mig inte att göra det här.
Ställ inte till en scen.
Se inte så chockad ut.
Låt inte Tom se dig.
Låt inte Tom se er.
Släpp mig inte.
Släpp inte taget om mig.
Gå inte.
Avbryt inte Tom.
Gå inte ut på framsidan.
Ge mig inte den där blicken.
Bli inte paranoid.
Lova att du inte blir arg.
Glöm inte din väska.
Glöm inte att använda tandtråd.
Smickra inte dig själv.
Drick inte det där.
Gör inte det här.
Gör inte detta.
Gör det inte.
Dö inte.
Var inte så negativ.
Var inte så negativa.
Var inte så lat.
Var inte så dramatisk.
Var inte oförskämd.
Var inte ohövlig.
Var inte ohyfsad.
Bli inte sårad. Tom är så där med alla.
Bli inte stött. Tom är så där med alla.
Var inte elak.
Var inte arg på mig.
Var inte fräck emot mig.
Var inte ohyfsad.
Spela inte förvånad.
Hälsa Tom att jag är färdig.
Säg till Tom att jag är färdig.
Säg till Tom att jag älskar honom.
Berätta för Tom att jag älskar honom.
Säg att du skämtar!
Berätta vad du såg.
Säg mig vad du tycker.
Berätta för mig om Tom.
Säg åt Mary att jag älskar henne.
Ta Tom till stationen.
Ta ut soporna.
Ta väl hand om Tom.
Ta hand om Tom.
Stanna bilen.
Sluta med det där.
Sluta upp med det där.
Sluta prata med mig.
Stanna, annars skjuter jag.
Sluta trakassera mig.
Sluta besvära mig.
Sluta kalla mig för Tom.
Sluta vara så dramatisk.
Sluta plåga mig.
Sluta tjata på mig.
Stanna här med Tom.
Underteckna på den här raden.
Signera på raden här.
Spela den sången igen.
Ryck upp dig.
Låt mig tänka en minut.
Låt mig fundera en minut.
Låt mig ta en titt.
Får jag se den där listan.
Låt mig hjälpa till.
Låt mig hjälpa dig upp.
Låt mig ta hand om Tom, okej?
Låt mig ringa min advokat.
Håll Tom utanför detta.
Håll Tom utanför det här.
Lämna min familj ifred.
Sänk rösten.
Håll dina händer borta från mig.
Ur vägen för mig.
Håll dig ur min väg.
Håll er ur min väg.
Släng iväg den bara.
Kasta den bara.
Ta bara ett djupt andetag.
Kom ned från scenen bara.
Följ bara mitt exempel.
Berätta bara inte för Tom.
Blunda bara.
Bromsa.
Gå och vänta i bilen.
Gå hem. Vila upp dig.
Gå och hämta lite handdukar.
Återgå till arbetet.
Få bort Tom härifrån.
Tar du dörren?
Sov lite.
Ta reda på vem Tom har pratat med.
Ta reda på var Tom är.
Ta reda på vad Tom vill.
Fyll i den här, tack.
Fyll i denna, tack.
Gör det snabbt.
Gör det fort.
Lugna dig.
Kom och träffa några av dina nya klasskamrater.
Kom och träffa allihop.
Kom tillbaka hit.
Ring mig när det är färdigt.
Ta det lugnt.
Jag bor inte i Finland.
Hon var inte snabb nog.
Hon var inte tillräckligt snabb.
Hans föräldrar älskar mig.
"Kunde du hämta en kopp kaffe åt mig?" "Visst. Så gärna."
Tom skrek åt Mary.
Tom skrek på Mary.
Tom kommer inte att stanna.
Tom lyssnar inte.
Tom kommer att bli överlycklig.
Tom kommer att vara här.
Tom var väldigt modig.
Tom hade rätt.
Tom var min hjälte.
Tom var gift på den tiden.
Tom var otrolig.
Tom var ofattbar.
Tom var fantastisk.
Tom avrättades i elektriska stolen.
Tom gavs en dödande elektrisk stöt.
Tom var deprimerad.
Tom är för tidigt född.
Tom blev arresterad.
Tom blev kidnappad.
Tom blev bortförd.
Tom blev bortrövad.
Tom vill leka.
Tom vill spela.
Tom vill ha hjälp.
Tom vill ha en kyss.
Tom vill ha en puss.
Tom ville träffa Mary.
Tom bleknade.
Tom blev blek.
Tom snavade och föll.
Tom försökte behålla lugnet.
Tom försökte rädda mig.
Tom försökte döda mig.
Tom tog av sig skjortan.
Tom tog av sig tröjan.
Tom stal dina pengar.
Tom stal era pengar.
Tom började skratta.
Tom låter utmattad.
Tom halkade och föll.
Tom borde ha varit här vid det här laget.
Tom borde vara här.
Tom sköt mig i benet.
Tom skakade på huvudet.
Tom skickade mig ett meddelande.
Tom verkar stressad.
Tom verkar trevlig.
Tom verkade trevlig.
Tom verkade borta.
Tom verkade vilse.
Tom såg videon.
Tom satt på trottoarkanten.
Tom rullade med ögonen.
Tom himlade med ögonen.
Tom lurade mig.
Tom lade ned boken.
Tom la ner boken.
Tom lovade att hjälpa.
Tom tog upp telefonen.
Tom tuppade av.
Tom svimmade.
Tom kolade av.
Tom dog.
Tom öppnade dörren.
Tom öppnade sin resväska.
Tom lyssnar aldrig på mig.
Tom hade aldrig en chans.
Tom hade aldrig någon chans.
Tom kom aldrig tillbaka.
Tom behöver vinna tid.
Tom behöver mig.
Tom behöver hjälp.
Tom behöver en tjänst.
Tom behövde pengar.
Tom behövde kontanter.
Tom måste stoppas.
Tom måste hjälpas.
Tom måste få hjälp.
Tom saknar dig.
Tom saknar Mary.
Tom har kanske rätt.
Tom fick mig att göra det.
Tom fick Mary att sluta.
Tom valde.
Tom gjorde sitt val.
Tom tog ett beslut.
Tom fattade ett beslut.
Tom sänkte rösten.
Tom ser sjuk ut.
Tom ser illamående ut.
Tom ser lättad ut.
Tom ser ut som du.
Tom ser skyldig ut.
Tom ser frustrerad ut.
Tom ser bekant ut.
Tom ser utmattad ut.
Tom ser utpumpad ut.
Tom ser slut ut.
Tom ser äcklad ut.
Tom ser annorlunda ut.
Tom ser förkrossad ut.
Tom såg förbryllad ut.
Tom ser förvirrad ut.
Tom ser konfys ut.
Tom ser konfunderad ut.
Tom ser omtumlad ut.
Tom ser irriterad ut.
Tom ser besvärad ut.
Tom ser arg ut.
Tom ser orolig ut.
Tom ser upphetsad ut.
Tom ser upprörd ut.
Tom ser lättad ut.
Tom såg bra ut.
Tom tittade på golvet.
Tom tittade i golvet.
Tom tittade på klockan.
Tom kollade på klockan.
Tom tittade på Mary.
Tom tittade på sin klocka.
Tom kollade på sin klocka.
Tom lånade mig den där DVD:n.
Tom bor på en båt.
Tom gillar det hett.
Tom gillar det varmt.
Tom gillar den varm.
Tom gillar det kallt.
Tom gillade den idén.
Tom tyckte om den idén.
Tom ljög för dig.
Tom släppte in mig.
Tom lämnade ett meddelande.
Tom lever ett stillsamt liv.
Tom vet var Mary är.
Tom vet att han har rätt.
Tom var medveten om riskerna.
Tom visste att jag var på väg.
Tom sparkade omkull en stol.
Tom behöll min tändare.
Tom gick just in.
Tom gick precis in.
Tom gick bara in.
Tom stirrade bara på Mary.
Tom dök precis upp.
Tom dök bara upp.
Tom försvann just.
Tom försvann bara.
Tom försvann precis.
Tom sitter inte i fängelse.
Tom är inte i häkte.
Tom sitter inte i häkte.
Det är inte Tom som bestämmer.
Tom är inte glad.
Tom är inte död.
Tom andas inte.
Tom är inte rädd för dig.
Tom är ingen främling.
Tom arbetar.
Tom är klarvaken.
Tom väntar på dig.
Tom väntar på er.
Tom väntar på Mary.
Tom är på övervåningen.
Tom har någonting på gång.
Tom är omöjlig att hindra.
Tom är omöjlig att stoppa.
Tom är ohejdbar.
Tom är för ung.
Tom är för långt borta.
Tom är deras ledare.
Det är Tom som bestämmer.
Tom är chef.
Tom är fortfarande skeptisk.
Tom gråter fortfarande.
Tom sover fortfarande.
Tom är fortfarande vid liv.
Tom är rädd.
Tom är precis här.
Tom är här.
Tom är mycket fotogenisk.
Tom har timlön.
Tom är på lastkajen.
Tom är på lastningsplatsen.
Tom är på väg hit.
Tom kommer inte.
Tom är inte rolig.
Tom har aldrig fel.
Tom är min make.
Tom är min man.
Tom är min hjälte.
Tom saknas.
Tom saknar ett finger.
Tom är eländig.
Tom är olycklig.
Tom är förtvivlad.
Tom är gift.
Tom tittar på mig.
Tom tittar på den.
Tom är bara rädd.
Tom är illa ute.
Tom är i knipa.
Tom har problem.
Tom är i duschen.
Tom är på sjukhuset.
Tom är uppe på vinden.
Tom ligger i koma.
Tom ignorerar dig.
Tom håller i en kniv.
Tom döljer någonting.
Tom kommer att klara sig.
Tom är rasande.
Tom är ursinnig.
Tom är mållös.
Tom är häpen.
Tom är förbluffad.
Tom är förstummad.
Tom är besviken.
Tom är desperat.
Tom är död.
Tom kommer tillbaka.
Tom är bakom dig.
Tom är knappt vid liv.
Tom är tillbaka i stan.
Tom är vid dörren.
Tom är på baren.
Tom är på flygplatsen.
Tom är föräldralös.
Tom är ett föräldralöst barn.
Tom är en gammal vän.
Tom är redan där.
Tom ska precis gå.
Tom är en smart grabb.
Tom är en stamkund.
Tom är en stamgäst.
Tom är fast anställd.
Tom är en bra grabb.
Tom är en bra vän.
Tom är miljardär.
Tom lade på telefonen.
Tom la på telefonen.
Tom la på i örat på Mary.
Tom hjälpte oss mycket.
Tom hjälpte mycket.
Tom höll Mary tätt.
Tom satte av mot dörren.
Tom hatar dig.
Tom hatar mig.
Tom har åkt fast för rattfylleri två gånger.
Tom måste gå hem.
Tom har svimmat.
Tom har tuppat av.
Tom har kolat av.
Tom har aldrig haft ett jobb.
Tom är skadad.
Tom har blivit skadad.
Tom gav Mary en kopp.
Tom hade inget val.
Tom högg tag i sin väska.
Tom grep tag i sin väska.
Tom ryckte till sig sin väska.
Tom hoppade av sin häst.
Tom satte sig i bilen.
Tom bor inte här.
Tom låter inte Mary gå och shoppa ensam.
Tom vet inte.
Tom har inget hem.
Tom hatar dig inte.
Tom hatar er inte.
Tom hatar inte dig.
Tom hatar inte er.
Tom dog ensam.
Tom berättade inte det för mig.
Tom såg det inte.
Tom såg inte det.
Tom nämnde inte det.
Tom nämnde inte Mary.
Tom dödade inte Mary.
Tom begick inte självmord.
Tom tog inte självmord.
Tom dödade ingen.
Tom dödade inte någon.
Tom gjorde det, eller hur?
Tom klappade ihop.
Tom tog knäcken på sig.
Tom kunde inte hitta Mary.
Tom kunde inte finna Mary.
Tom skulle kunna vara var som helst.
Tom skulle kunna vara en polis.
Tom kollade tiden.
Tom sprang efter Mary.
Tom kan inte gå.
Tom kan inte stanna.
Tom kan inte se dig.
Tom får inte se dig.
Tom kan inte träffa dig.
Tom får inte träffa dig.
Tom kan inte skada dig.
Tom kan inte skada mig.
Tom får inte skada mig.
Tom hör dig inte.
Tom kan inte höra dig.
Tom kan inte vara allvarlig.
Tom kan inte vara seriös.
Tom kan visa dig runt.
Tom kan höra dig.
Tom kan höra er.
Tom kom för att hjälpa.
Tom frågade ut mig.
Hajar är goda simmare.
Jag vill inte vara rik.
Du har många vänner.
Mary har många vänner.
Ring dem i kväll.
Det är nästan omöjligt.
Det är närapå omöjligt.
Tom sa att han inte var intresserad av Mary, men det verkade som att han alltid tittade åt den del av rummet som hon var i.
Detta är inkorrekt.
Det här är inkorrekt.
Detta är oriktigt.
Det här är oriktigt.
Detta är felaktigt.
Det här är felaktigt.
Det här är inte rätt.
Det här är inte korrekt.
Det här är inte riktigt.
Det här är inte rätt.
Detta är inte rätt.
Detta stämmer inte.
Det här stämmer inte.
Tom kommer inte att döda någon annan.
Varför svarar du inte?
Var finns närmaste hotell?
Jag är trött eftersom jag arbetade för mycket.
Detta är skandalöst!
Det här är skandalöst!
Han berättade aldrig för någon.
Jag lovar. Jag kommer aldrig att göra det igen.
Tom är fortfarande vaken.
Tom är fortfarande uppe.
Tom är fortfarande vaken.
Jag älskar det norska språket!
Jag älskar det norska språket!
Det är min fru.
Jag är redan sen.
Jag vet var han är.
Var täckte du över dom?
Han är irriterande.
Han är besvärlig.
Hon gjorde så gott hon kunde.
Han deltog i en nätundersökning.
Hur mår din patient?
Hur är det med Tom?
Hur går det för Tom?
Hur går det med skolan?
Hur går det på skolan?
Hur går det i skolan?
Hur går det?
Hur mår du?
Hur känner du dig?
Hur kom du hit?
Hur tog du dig hit?
Hur skulle du veta?
Hur mycket kostar det där?
Hur mycket är det där?
Hur mycket vill du ha?
Hur mycket vill ni ha?
Hur mycket kostade det?
Hur mycket kostade den där?
Hur många tog du?
Hur många fick du?
Hur många fick du tag på?
Hur länge var Tom här?
Hur länge har vi på oss?
Hur lång tid har vi?
Hur lång tid har vi på oss?
Hur lång tid har du på dig?
Hur länge har vi på oss?
Hur lång tid har vi?
Hur är detta relevant?
Hur är det relevant?
Hur svårt kan det vara?
Hur ser det här ut?
Hur känns det?
Hur känns det där?
Hur fungerar det?
Hur ser det ut?
Hur tror du att jag känner?
Hur tror ni att jag känner?
Hur tror du att jag känner mig?
Hur tror ni att jag känner mig?
Hur känner du Tom?
Hur känner ni Tom?
Hur visste du?
Hur gissade du?
Hur kunde du gissa?
Hur fick du tag på dem där?
Hur kom du in hit?
Hur kom ni in hit?
Hur tog du dig in hit?
Hur tog ni er in hit?
Hur hittade ni oss?
Hur hittade du oss?
Hur hittade du Tom?
Hur hamnade du här?
Hur hamnade ni här?
Hur träffade Tom Mary?
Hur såg Tom ut?
Hur visste Tom det?
Hur hittade Tom oss?
Hur fick Tom reda på det?
Hur hände det där?
Hur löste sig allt?
Hur gick det med allt?
Hur gjorde du det?
Hur gjorde ni det?
Hur vet du det?
Hur vet ni det?
Hur kan vi tacka er?
Hur kan vi tacka dig?
Hur kan vi rädda Tom?
Hur kan vi göra det?
Hur kan detta vara sant?
Hur kan det vara sant?
Hur kan jag hjälpa till?
Hur kan jag hjälpa?
Hur illa var det?
Hur dåligt var det?
Hur illa är det?
Hur mår du nu?
Har du sovit?
Har du sett Tom?
Har du sett Tom än?
Har ni sett Tom än?
Har du sett det här?
Har du hört från Tom?
Har ni hört från Tom?
Har du hittat någonting?
Har ni hittat någonting?
Har du varit i Boston?
Har ni varit i Boston?
Har du rökt?
Har Tom blivit skadad?
Har Tom skadats?
Vill du inte åka?
Känner du inte igen Tom?
Känner ni inte igen Tom?
Tycker du inte om mig?
Vet du inte vem jag är?
Vet ni inte vem jag är?
Bryr du dig inte?
Ser Tom förvirrad ut?
Vet Tom?
Vet Tom om det?
Vet Tom än?
Vet Tom vem jag är?
Blir du ledsen av det?
Gör det dig ledsen?
Gör det er ledsna?
Blir ni ledsna av det?
Spelar det verkligen någon roll?
Spelar det någon roll?
Vill du hänga?
Vill ni hänga?
Vill du ha barn?
Vill du ha ett jobb?
Vill du ha ett arbete?
Ser du någonting?
Ser ni någonting?
Lovar du?
Lovar ni?
Äger du ett handeldvapen?
Äger du ett eldhandvapen?
Behöver du någonting?
Behöver ni någonting?
Behöver du en hand?
Saknar du Tom?
Saknar ni Tom?
Älskar du Tom?
Älskar ni Tom?
Gillar du Tom?
Tycker du om Tom?
Tycker du om robotar?
Vet du vem han var?
Vet ni vem han var?
Känner du Tom?
Känner du till Tom?
Måste du gå nu?
Måste ni gå nu?
Måste ni åka nu?
Måste du åka nu?
Har du några vapen?
Har du några kontanter?
Har du en telefon?
Har ni en telefon?
Tvivlar du på mig?
Använder du droger?
Klandrar du Tom?
Förebrår du Tom?
Lägger du skulden på Tom?
Tror du på mig nu?
Tror ni på mig nu?
Behöver vi en plan B?
Känner vi dig?
Känner vi er?
Har vi något val?
Ser jag OK ut?
Ser jag bra ut?
Måste jag betala dig?
Måste jag betala er?
Vann du trofén?
Vann du kapplöpningen?
Vann du kappkörningen?
Varnade du Tom?
Provade du det?
Berättade du för Tom?
Såg du Tom?
Träffade du Tom?
Har du gått ned i vikt?
Kände du Tom?
Kände du Tom väl?
Kände ni Tom väl?
Kysste du Mary?
Pussade du Mary?
Dödade du Tom?
Hörde du det?
Hade du roligt?
Hade du kul?
Fick du checken?
Fick ni checken?
Fattade du?
Hittade du din handväska?
Hittade du din börs?
Hittade du Tom?
Ringde du någonsin Tom?
Gjorde du det här?
Var det du som gjorde det här?
Köpte du Tom en hund?
Köpte ni Tom en hund?
Köpte du en hund till Tom?
Köpte ni en hund till Tom?
Köpte du en nya bil?
Köpte ni en ny bil?
Såg du den på riktigt?
Såg du det på riktigt?
Hotade Tom dig?
Såg Tom dig?
Sa Tom varför?
Blev Tom skadad?
Skadades Tom?
Förlät Tom dig?
Sa Tom det?
Kom Tom tillbaka?
Ringde Tom?
Har Tom ringt?
Sa de varför?
Sa de när?
Sa de hur?
Hittade dom någonting?
Hittade de någonting?
Skadades någon?
Gick det bra i dag?
Skrev jag det där?
Missade jag någonting?
Missade jag mycket?
Gjorde jag det där?
Var det jag som gjorde det där?
Berättade någon för Tom?
Sa någon någonting?
Skadades någon?
Gjorde någon sig illa?
Skulle jag kunna få en servett?
Kan du vakta ungarna?
Kan du passa barnen?
Kan ni passa barnen?
Kan du se dem?
Kan ni se dem?
Kan du laga en toalett?
Kan du ta reda på det?
Kan vi bara gå hem?
Har vi råd med det nu?
Kan Tom hjälpa oss?
Kan Tom få en hund?
Kan jag tänka på det?
Kan jag tänka på saken?
Kan jag få prata med dig?
Kan jag sitta ned?
Kan jag komma med dig?
Kan jag hämta er någonting?
Kan jag hämta dig någonting?
Kan jag få en hund?
Kan jag ringa upp dig?
Kan någon verifiera det?
Kan någon intyga det?
Kan något bekräfta det?
Kan någon bestyrka det?
Kan någon bevisa det?
Kan någon bevisa riktigheten av det?
Hotar du mig?
Hotar ni mig?
Jobbar du fortfarande med Tom?
Arbetar du fortfarande med Tom?
Är du fortfarande gift?
Är ni fortfarande gifta?
Är du fortfarande arg på mig?
Är ni fortfarande arga på mig?
Är du fortfarande hemma?
Är ni fortfarande hemma?
Är du hungrig över huvud taget?
Stöter du på mig?
Ska du ut?
Är du rädd än?
Är ni rädda än?
Följer du efter mig?
Följer ni efter mig?
Väntar du på Tom?
Gråter du?
Grinar du?
Kommer ni med oss?
Kommer du med oss?
Kommer du eller inte?
Rodnar du?
Är du en idiot?
Är du rädd för mig?
Är du polis?
Är du polisman?
Ska vi åka långt?
Ska vi gå långt?
Är vi vänner?
Är vi färdiga här?
Är det där mina örhängen?
Är de där till mig?
Är de där för mig?
Är de där åt mig?
Tydligen är jag adopterad.
Talar jag för snabbt?
Pratar jag för snabbt?
Kommer jag att dö?
Stör jag dig?
Stör jag er?
Stör jag dig?
Skulle Tom gilla det?
Skulle Tom tycka om det?
Varför frågar du det?
Varför skulle du fråga det?
Varför skulle Tom hjälpa oss?
Varför åker inte Tom?
Varför ger sig Tom inte iväg?
Varför ge dem någonting?
Jag kan väl skjutsa dig?
Varför skjutsar inte jag dig?
Varför sa Tom det?
Varför sa Tom så?
Varför är du hemma?
Varför är ni hemma?
Vems sida är du på?
På vems sida är du?
På vems sida är ni?
Vems sida är ni på?
Vems telefon är det där?
Vems idé var det?
Vems är de?
Vem är den här killen?
Vem är redo att beställa?
Vem håller utkik?
Vem är på vakt?
Vem går på vakt?
Vem skulle bry sig?
Var är väskan?
Var är mitt te?
Var är min telefon?
Var är min golfbag?
Var är min bil?
Var är alla?
Var är allihopa?
Var är allesammans?
Var ska jag lägga den?
Var bodde du?
Var bodde ni?
Var växte du upp?
Var växte ni upp?
Var fick du tag på den där?
Var hittade du Tom?
Var fann du Tom?
Vart gick Tom?
Var kom den ifrån?
Var kom det ifrån?
Var kan jag hitta Tom?
Vart är du på väg?
Var är vi nu?
Var är Toms saker?
Var är de?
Var är bilnycklarna?
Var är mina saker?
När är begravningen?
När var det?
När kommer Tom?
När behöver Tom den?
När behöver Tom det?
När börjar vi?
När startar vi?
När sa du det?
När sa ni det?
När sa du det där?
När sa ni det där?
När fick du den här?
När fick ni den här?
När frågade du Tom?
När sa Tom det?
När rymde Tom?
Vad har du?
Vad har du gjort?
Vad har ni gjort?
Vad är din plan?
Vad är er plan?
Vad hette du nu igen?
Vad var det du heter nu igen?
Vad är det för fel med det?
Vad är det med Tom?
Vad är Toms problem?
Vad heter Tom i efternamn?
Varför gömmer sig Tom?
Vad är det Tom gömmer sig för?
Vad har Tom hittat?
Vad gör Tom här?
Vad är den här till?
Vad används den här till?
Vadan denna panik?
Vad är avbrottet?
Vad är alternativet?
Vad är det som luktar?
Vad är det där för lukt?
Var har du fått det där ärret ifrån?
Var kommer det där ärret ifrån?
Vad är det som tar så lång tid?
Vad är det som tar en sådan tid?
Vad är det som är så kul?
Vad är det som är så roligt?
Vad är min belöning?
Varför dröjer Tom?
Vad uppehåller Tom?
Hur är den?
Hurdan är den?
Hur ser den ut?
Hur är det?
Hur känns det?
Vad handlar det om?
Vad finns där inne?
Vad finns på insidan?
Vad heter han?
Vad är du bra på?
Vi ska vi göra?
Vad ska vi ta oss till?
Vad var Toms plan?
Vad var problemet?
Vad fanns inuti?
Vad skrämde dig?
Vad dödade Tom?
Vad var det som Tom dödade?
Vad är det här för?
Vad är det här till?
Vad är detta för?
Vad är detta till?
Vad är det som pågår här?
Vad är allt det här?
Vad är allt detta?
Vad har du hört?
Vad händer i morgon?
Vad hände sen?
Vilken årskurs är Tom i?
Exakt vad är det där?
Vad mer behöver du?
Vad mer sa Tom?
Vad mer kan du göra?
Vad mer kan ni göra?
Vad minns du?
Vad minns ni?
Vad behöver du veta?
Vad vet du?
Vad har vi här?
Vad gör vi nu?
Vad är jag skyldig dig?
Vad är jag skyldig er?
Vad gör jag härnäst?
Vad gör jag sen?
Vad bryr jag mig om det?
Vad såg du?
Vad lärde du dig?
Vad träffade du?
Vad kallade du mig?
Vad kallade ni mig?
Vad missade vi?
Vad ville Tom?
Vad ville Tom ha?
Vad sa Tom?
Vad visste Tom?
Vad gjorde Tom?
Vad ville de?
Vad har vi för val?
Vad kan du ge mig?
Vad för dig hit?
Vad skriver du?
Vad har du på dig?
Vad har du på dig för kläder?
Vad är du rädd för?
Vad är ni rädda för?
Vad gör vi?
Vad är de där?
Stod ni två nära varandra?
Blev du beskjuten?
Blev Tom mördad?
Var Tom ensam?
Blev någon dödad?
Så vad hände?
Så vad gjorde du?
Borde inte du gå hem?
Borde inte ni gå hem?
Borde inte du åka hem?
Borde inte ni åka hem?
Ska vi beställa?
Är inte det planen?
Är det inte det som är planen?
Är det där Tom?
Kan de se oss?
Du skulle ha sett henne.
Jag ringde i förväg.
Jag kan knappt andas.
Jag kan höra vinden.
Jag kan hjälpa dig.
Jag kan inte tillåta det.
Jag kan inte svara på det.
Jag kan inte vara säker.
Jag kan inte göra mer.
Jag kan inte göra det själv.
Jag klarar det inte själv.
Jag kan inte göra det här längre.
Jag kan inte göra detta.
Jag kan inte göra det här.
Jag kan inte rita en fågel.
Jag kan inte hitta den.
Jag kan inte hitta det.
Jag kan inte bli inblandad.
Jag hör ingenting.
Jag kan inte höra någonting.
Jag kan inte behålla det här.
Jag kan inte behålla den här.
Jag kan inte leva med det.
Jag hinner inte.
Jag dubbelkollade det.
Jag kollade det två gånger.
Jag kontrollerade det två gånger.
Jag kommer hit varje dag.
Jag skulle kunna kyssa dig.
Jag kunde inte bry mig mindre.
Jag skulle inte kunna bry mig mindre.
Det rör mig inte i ryggen.
Jag kunde inte ljuga för dig.
Jag kunde inte ljuga för er.
Jag kunde inte säga nej.
Jag kan inte se någonting.
Jag kunde inte se någonting alls.
Jag kunde inte stå.
Jag gjorde ingenting.
Jag gjorde dig en tjänst.
Jag bad inte om detta.
Jag bad inte om det här.
Jag gjorde det inte.
Jag behövde inte gå.
Jag behövde inte åka.
Jag var inte tvungen att gå.
Jag var inte tvungen att åka.
Jag dödade inte någon.
Jag dödade inte Tom.
Jag menade inte något av det.
Jag flyttade inte på någonting.
Jag behövde inte din hjälp.
Jag behövde inte er hjälp.
Jag sa inget.
Jag sa ingenting.
Jag sov inte bra.
Jag rörde inte Tom.
Jag ville inte ha mjölk.
Jag skrev ingenting.
Jag skrev inte någonting.
Jag gör det hela tiden.
Jag tror inte på det.
Jag förtjänar inte detta.
Jag förtjänar inte det här.
Jag känner mig inte sjuk.
Jag känner mig inte särskilt lycklig.
Jag får inte så mycket post.
Jag måste inte vara här.
Jag känner inte Tom.
Jag vet inte vad ni vill att jag ska säga.
Jag vet inte vad du vill att jag ska säga.
Jag har inget emot att hjälpa till.
Jag behöver ingen hjälp.
Jag känner inte igen det.
Jag känner inte igen den.
Jag litar inte på någon.
Jag vill inte ha det här.
Jag vill inte ha den här.
Jag vill inte ha denna.
Jag vill inte ha detta.
Jag kör en hybrid.
Jag kör en hybridbil.
Jag känner mig illamående.
Jag kände mig skyldig.
Jag konstaterade en sak.
Jag fick reda på någonting.
Jag kom underfund med någonting.
Jag hittade din dagbok.
Jag fann din dagbok.
Jag gav Tom ett val.
Jag gav inte Tom något val.
Jag blev betalad i dag.
Jag antar att Tom inte är hemma.
Jag antar att du har rätt.
Jag var tvungen att göra någonting.
Jag hatar att vara dum.
Jag hatar min röst.
Jag hatar folk som Tom.
Jag hatar människor som Tom.
Jag hatar personer som Tom.
Jag hatar överraskningar.
Jag har ett tillkännagivande.
Jag har en kungörelse.
Jag har ett meddelande.
Jag har en annan idé.
Jag har en till fråga.
Jag har en annan fråga.
Jag har ryggproblem.
Jag har massor med vänner.
Jag har min egen teori.
Jag har så många idéer.
Jag måste ändra på mig.
Jag måste göra det själv.
Jag måste göra det här själv.
Jag måste göra detta själv.
Jag måste åka hem.
Jag måste ta mig hem.
Jag måste gå.
Jag måste få träffa Tom.
Jag måste träffa Tom.
Jag har arbete att göra.
Jag hör skratt.
Jag hörde ett ljud.
Jag hörde ett oljud.
Jag hörde det på tv.
Jag hörde meddelandet.
Jag hörde röster.
Jag hoppas att det inte är sant.
Jag hoppas att det där inte är sant.
Jag hoppas att Tom är okej.
Jag hoppas att Tom säger ja.
Jag hoppas att vi hittar Tom.
Jag hoppas att vi finner Tom.
Jag hoppas att du är hungrig.
Jag hoppas att du har rätt.
Jag lånade den precis.
Jag lånade den bara.
Jag lånade den just.
Jag kan bara inte sova.
Jag kan inte sova bara.
Jag kunde bara inte säga nej.
Jag vet bara inte.
Jag hittade den precis.
Jag hittade det just.
Jag hittade den just.
Jag hittade det precis.
Jag fick precis sparken.
Jag fick precis ditt mejl.
Jag fick precis ditt mail.
Jag tjänade precis tre lax.
Jag träffade honom precis.
Jag behöver bara en minut.
Jag behöver bara hitta Tom.
Jag öppnade den precis.
Jag stötte precis min tå.
Jag stötte precis tån.
Jag vill bara gå hem.
Jag vill bara åka hem.
Jag vill bara vila.
Jag vill bara prata.
Jag ville bara ha pengar.
Jag visste att jag inte var galen.
Jag visste vad du menade.
Jag visste vad ni menade.
Jag visste att du skulle bli arg.
Jag visste att du skulle gilla det.
Jag visste att du skulle gilla den.
Jag visste att du skulle tycka om det.
Jag visste att du skulle tycka om den.
Jag kände din far.
Jag kände din fader.
Jag kände din pappa.
Jag vet allt om dig.
Jag vet allting om dig.
Jag kan allt det här.
Jag vet allt det här.
Jag kan allt detta.
Jag vet allt detta.
Jag vet hur gammal Tom är.
Jag vet hur detta fungerar.
Jag vet hur det här funkar.
Jag vet att det här är svårt.
Jag vet att detta är svårt.
Jag vet att det är svårt.
Jag känner Tom personligen.
Jag vet vad jag vill.
Jag vet vad jag vill ha.
Jag vet vad som dödade Tom.
Jag vet vad som är rätt.
Jag vet vad som är fel.
Jag vet vem som gjorde det.
Jag vet att du mår dåligt.
Jag vet att du är upptagen.
Jag vet att ni är upptagna.
Jag vet att du har rätt.
Jag vet att du är upprörd.
Jag vet att ni är upprörda.
Jag lämnade dig ett meddelande.
Jag gillar att vara upptagen.
Jag gillar hur Tom tänker.
Jag tycker om hur Tom tänker.
Jag gillar den där tröjan.
Jag gillar den där skjortan.
Jag gillar att vara förberedd.
Jag gillar din hund.
Jag tycker om din hund.
Jag gillar ditt hår.
Jag gillar din hatt.
Jag tycker om din hatt.
Jag gillar din scarf.
Jag gillar din halsduk.
Jag gillar din sjal.
Jag gillar din sjalett.
Jag tycker om din scarf.
Jag tycker om din halsduk.
Jag tycker om din sjal.
Jag tycker om din sjalett.
Jag gillade den där filmen.
Jag gillade den filmen.
Jag gillade din historia.
Jag tyckte om din historia.
Jag låste dörren på framsidan.
Jag tappade ett örhänge.
Jag tappade tidsuppfattningen.
Jag älskar utmaningar.
Jag älskar Mary så mycket.
Jag älskar den där klänningen.
Jag älskar den filmen.
Jag älskar den scarfen.
Jag älskar den halsduken.
Jag älskar den sjalen.
Jag älskar den sjaletten.
Jag älskar den sången.
Jag älskar den berättelsen.
Jag älskar den historian.
Jag älskar den sagan.
Jag älskar det här jobbet.
Jag älskar detta jobb.
Jag älskar detta arbete.
Jag älskar det här arbetet.
Jag älskar den här delen.
Jag älskar denna del.
Jag älskar den här staden.
Jag älskar denna stad.
Jag älskar er båda.
Jag älskar dina ögon.
Jag älskar ditt hår.
Jag gjorde några ändringar.
Jag gjorde den där.
Jag kanske kommer att prata med Tom.
Jag kanske pratar med Tom.
Jag saknar Tom så mycket.
Jag saknar dig, Tom.
Jag behöver en advokat.
Jag behöver en huvudvärkstablett.
Jag behöver min jacka.
Jag behöver min rock.
Jag behöver min kappa.
Jag behöver lite sömn.
Jag behöver lite vatten.
Jag behöver bilnycklarna.
Jag behöver få träffa Tom.
Jag behöver träffa Tom.
Jag behöver dig här.
Jag behöver att du går hem.
Jag såg dig aldrig.
Jag såg aldrig dig.
Jag såg aldrig er.
Jag såg er aldrig.
Jag tar aldrig sovmorgon.
Jag rörde den aldrig.
Jag rörde aldrig Tom.
Jag gick aldrig och la mig.
Jag gick aldrig och lade mig.
Jag föredrar att gå.
Jag läste din rapport.
Jag behöver verkligen din hjälp.
Jag behöver verkligen er hjälp.
Jag sa stick.
Jag räddade ditt liv.
Jag såg allt.
Jag såg Tom i dag.
Jag träffade Tom i dag.
Jag träffade Tom i kväll.
Jag såg Tom i kväll.
Jag såg vad Tom gjorde.
Jag såg vad du gjorde.
Jag förstår vad problemet är.
Jag träffar Tom varje dag.
Jag ser Tom varje dag.
Jag skickade iväg Tom.
Jag skickade hem Tom.
Jag borde vila upp mig lite.
Jag borde vila mig lite.
Jag borde få mig lite vila.
Jag borde inte vara här.
Jag gillar det fortfarande inte.
Jag tycker fortfarande inte om det.
Jag stal den från Tom.
Jag stal det från Tom.
Jag sträckte ut armarna.
Jag sträckte ut benen.
Jag pratade med Tom.
Jag talade med Tom.
Jag berättar allt för Tom.
Jag tror att jag gillar dig.
Jag tror att jag är förälskad.
Jag tror att jag är kär.
Jag tror att Mary tycker om mig.
Jag tror att Mary gillar mig.
Jag tror att Tom ljuger.
Jag tror att Tom gick.
Jag tror att Tom ljög för oss.
Jag tycker vi borde göra mer än så.
Jag tror att vi borde gå.
Jag tror att vi borde åka.
Jag tror att det är bäst att du går.
Jag tycker att du är trevlig.
Jag tycker att du är snäll.
Jag tyckte att det var gott.
Jag tyckte att det var bra.
Jag trodde att du slutade.
Jag trodde att du slutat.
Jag trodde du var van vid att bo i husvagn.
Jag berättade sanningen för Tom.
Jag sa åt dig att gå.
Jag sa åt er att gå.
Jag sa åt dig att ge dig iväg.
Jag sa åt er att ge er iväg.
Jag tog Tom till sjukhuset.
Jag förstår helt och hållet.
Jag försökte varna dig.
Jag försökte varna er.
Jag vill ha en advokat.
Jag vill be om ursäkt.
Jag vill vara här.
Jag vill tro dig.
Jag vill tro er.
Jag vill komma hem.
Jag vill drömma.
Jag vill åka tillbaka.
Jag vill gå tillbaka.
Jag vill träffa Tom.
Jag vill träffa Tom.
Jag var ironisk.
Jag var artig.
Jag var hövlig.
Jag föddes här.
Jag var på området.
Jag tar den.
Jag skulle dö utan dig.
Jag skulle dö utan er.
Jag skulle hjälpa dig om jag kunde.
Jag skulle hjälpa er om jag kunde.
Jag skulle vilja tro dig.
Jag skulle vilja tro er.
Jag skulle vilja träffa Tom.
Jag skulle vilja se Tom.
Jag kommer att vara hos Tom.
Jag är hos Tom.
Jag klarar mig.
Jag kommer att vara här.
Jag är här.
Jag stannar här.
Jag är på mitt kontor.
Jag kommer att vara på mitt kontor.
Jag ringer efter en taxi åt dig.
Jag ringer en taxi åt dig.
Jag ska kolla igen.
Jag ska göra det nu.
Jag kommer att drömma om dig.
Jag ska hämta min jacka.
Jag ska ta min jacka.
Jag ska hämta min rock.
Jag ska ta min rock.
Jag ska hämta min kappa.
Jag ska ta min kappa.
Jag hämtar mina nycklar.
Jag hämtar nycklarna.
Jag ska hämta mina nycklar.
Jag ska hämta nycklarna.
Jag fixar en.
Jag hämtar en.
Jag hämtar lite is.
Jag hämtar boken.
Jag ska hämta boken.
Jag hämtar bilen.
Jag ska hämta bilen.
Jag går och frågar Tom.
Jag ska gå och fråga Tom.
Jag kommer att gå och fråga Tom.
Jag går först.
Jag kommer att gå först.
Jag ska gå och handla.
Jag ska gå och shoppa.
Jag följer med dig.
Jag kommer att följa med dig.
Jag ska följa med dig.
Jag ska ta hand om det.
Jag tar hand om det.
Jag tar hand om det här.
Jag kommer att ta hand om det här.
Jag ska ta hand om det här.
Jag kommer att hjälpa dig.
Jag håller dig informerad.
Jag håller dig à jour.
Jag undersöka det.
Jag forska i det.
Jag ska ringa några samtal.
Jag betalar det dubbla.
Jag betalar extra.
Jag ska betala extra.
Jag kommer att betala extra.
Jag betalar på mitt eget sätt.
Jag ska betala dig.
Jag hämtar upp Tom.
Jag kommer att hämta upp Tom.
Jag ska hämta upp Tom.
Jag ska skjuta dig.
Jag skjuter dig.
Jag kommer att skjuta dig.
Jag pratar med Tom.
Jag ska prata med Tom.
Jag kommer att prata med Tom.
Jag berättar för Tom senare.
Jag ska berätta för Tom senare.
Jag ska berätta för dig.
Jag kommer att berätta för dig.
Jag berättar för dig.
Jag väntar här.
Jag kommer att vänta här.
Jag ska jobba på det.
Jag är lite upptagen.
Jag är lite tidig.
Jag är musiker.
Jag är en tålmodig man.
Jag är fotograf.
Jag är socialarbetare.
Jag är alldeles ensam nu.
Jag är helt ensam nu.
Jag är redan rik.
Jag är oskyldig.
Jag är en oskyldig man.
Jag är hemskt trött.
Jag ringer polisen.
Jag kommer till dig.
Jag gör mina läxor.
Jag är lealös.
Jag är mjuk i lederna som en akrobat.
Jag väntar ett samtal.
Jag känner mig hungrig.
Jag är färdig.
Jag ska skaffa katt.
Jag håller på att bli bättre.
Jag är glad att vi är överens.
Jag är glad att du är här.
Jag håller på att bli galen.
Jag blir galen.
Jag ska gå nu.
Jag kommer att gå nu.
Jag går nu.
Jag ska försöka.
Jag kommer att försöka.
Jag följer med Tom.
Jag är så gott som aldrig hemma.
Jag är nästan aldrig hemma.
Jag är här varje kväll.
Jag är här för att be om ursäkt.
Jag är här för att hjälpa dig.
Jag är här för att hjälpa er.
Jag är på vinden.
Jag är på vindsvåningen.
Jag är bara en taxichaufför.
Jag är bara ärlig.
Jag chansar bara.
Jag är bara lat.
Jag är precis som du.
Jag är något av en ensamvarg.
Jag är sen till jobbet.
Jag är sen till arbetet.
Jag håller på att bli galen.
Jag är arg på dig.
Jag är ingen tiggare.
Jag ger inte upp.
Jag kommer inte att dö.
Jag ska inte dö.
Jag är precis här.
Jag är trött på det här.
Jag har fått nog av det här.
Jag är så generad.
Jag är så stolt över dig.
Jag är mördaren.
Jag har sett det här förut.
Jag har sett detta förut.
Toms farfar och Marys farfar slogs tillsammans i andra världskriget.
Toms farfar och Marys morfar slogs tillsammans i andra världskriget.
Toms morfar och Marys farfar slogs tillsammans i andra världskriget.
Toms morfar och Marys morfar slogs tillsammans i andra världskriget.
Vi är sena.
Jag är här.
Jag är precis här.
Vi är redo för detta.
Vi är i en konjunktursvacka.
Vi är i en recession.
Vi är i en lågkonjunktur.
Vi kommer att försöka.
Vi kommer att överleva.
Vi har pratat färdigt.
Vi kommer att vara där.
Vi klarar oss.
Vi kommer att klara oss.
Vi förstår.
Vi borde sätta upp en fälla.
Vi borde sätta igång.
Vi borde komma igång.
Vi borde ge oss av.
Vi borde ringa Tom.
Vi tummade på det.
Vi tog varandra i handen på det.
Vi måste prata med er om Tom.
Vi måste prata med dig om Tom.
Vi måste tala med er om Tom.
Vi måste tala med dig om Tom.
Vi måste skynda oss.
Vi måste hjälpa Tom.
Vi måste gå.
Vi måste göra det igen.
Vi matade just babyn.
Vi matade just barnet.
Vi måste flytta.
Vi måste förflytta oss.
Vi måste komma på ett sätt att få den här maskinen att fungera under vatten.
Vi måste göra bättre ifrån oss.
Vi har saker att göra.
Vi har inga hemligheter.
Vi har varit uppe hela natten.
Vi vill inte skrämma bort barnen.
Vi insåg inte att vi var så högljudda.
Det kan vi inte göra.
Vi kan göra det där.
Sedermera antog han en ny identitet.
Han har inte hatt på sig.
Jag vill bara ha roligt.
Jag vill bara ha kul.
Du är min enda glädje.
Låt oss göra affärer.
Det är inget problem.
Det är inga problem.
Du är konstig.
Du är en sådan flörtis.
Du kommer med undanflykter.
Du är så kinkig.
Du är så kräsen.
Du är så paranoid.
Ni är så paranoida.
Du kör så mycket med folk.
Du domderar så mycket.
Du är smartare än jag.
Du är smartare än jag.
Du är smartare än vad jag är.
Du har slut på ursäkter.
Ni har slut på ursäkter.
Du hjälper inte till.
Ni hjälper inte till.
Du är partisk.
Du babblar.
Du pladdrar.
Du är en snobb.
Du kommer att klara dig.
Du borde lita på mig.
Du ser så vacker ut.
Du måste lämna Boston.
Du skrämmer mig inte.
Ni skrämmer mig inte.
Du kan ta det.
Du kan ta den.
Vem som än använder den här tandborsten är inte min mor.
Det skulle kunna vara kul.
Det skulle kunna vara roligt.
Det känns riktigt bra.
Det var värt det.
Det är en plan.
Det där är ett gammalt skämt.
Det är okej.
Det är mycket.
Vad gjorde Tom med pengarna?
Vad gjorde Tom av pengarna?
De där är trevliga.
De där är fina.
Det här är konstigt.
Detta är konstigt.
Detta är underligt.
Det här är underligt.
Det här är väldigt färskt.
Det här är riktigt illa.
Detta är riktigt illa.
De kommer med undanflykter.
De slingrar sig.
De överstegrar.
De kör fast.
De är dyra.
Snälla kör in till trottoarkanten.
Mary kom självmant.
Mary kom själv.
Här kommer Tom.
Han slåss mot väderkvarnar.
Hon väntar.
Det varierar en hel del.
Det hände så fort.
Det hände så snabbt.
Ta bara en.
Du måste göra som jag säger.
Ni måste göra som jag säger.
Litar du på Tom?
Han föste iväg henne.
Det här är brevet från min vän.
Jag gjorde det frivilligt.
Det var ett insidejobb.
Det var ett internt jobb.
Var trevligare mot din syster.
Var trevligare mot er syster.
Ät dina grönsaker.
De andra barnen kallar henne Piggy.
De andra barnen kallar henne Nasse.
Lova mig att du inte berättar för henne.
Hon har ingen biljett.
Han har ingen biljett.
Hur ofta tvättar du dina jeans?
Han gillar indisk mat.
Var trevlig.
Mitt marsvin var min första flickvän.
Ser du porträttet?
En hunds nos är väldigt känslig.
Hon är en fanatiker.
Han kan tala med andar.
Han dricker inte.
Ett DNA-test visade att han var oskyldig.
Har du en kofot i verktygslådan?
Han håller på att bli skallig.
Det är dödligt gift!
Hur illa kan det vara?
Hur dåligt kan det vara?
Hur dålig kan den vara?
Han är inget helgon.
Jag fick ett F i kemi.
Jag fick C i engelska.
Jag fick B i fysik.
Jag fick A på min uppsats.
Jag uppskattar ditt jobb.
Jag uppskattar ditt arbete.
Jag uppskattar ert arbete.
Jag uppskattar din tid.
Jag uppskattar hjälpen.
Jag uppskattar det.
Jag har försökt att lösa det här problemet i timmar.
Försvinn från min gräsmatta!
Han är mörk och snygg.
Släpp henne.
Jag skulle vilja pröva det här.
Jag skulle vilja prata med Tom.
Jag skulle vilja tala med Tom.
Jag skulle vilja stå upp.
Jag skulle vilja träffa Tom nu.
Jag skulle vilja se det.
Jag skulle vilja följa med dig.
Jag skulle vilja hjälpa till.
Jag skulle vilja hjälpa dig.
Jag skulle vilja följa med Tom.
Jag skulle vilja gå hem nu.
Jag skulle vilja låna den här.
Jag skulle vilja låna detta.
Jag skulle vilja vara ensam.
Jag skulle vilja ställa dig några till frågor.
De hade inga skägg, inget hår och inga ögonbryn.
Jag trodde att Tom skulle sova över i Boston.
Jag trodde att Tom skulle stanna lite längre.
Jag trodde att Tom skulle tala bättre franska än Mary.
Jag trodde att Tom skulle sova till mitt på dagen.
Jag trodde att Tom skulle komma.
Jag trodde att Tom skulle dyka upp.
Jag trodde att Tom skulle säga det.
Jag trodde att Tom skulle säga hej.
Jag trodde att Tom skulle säga hej till Mary.
Jag trodde att Tom skulle komma ihåg.
Jag trodde att Tom skulle minnas.
Jag trodde att Tom skulle plantera de där blommorna nära eken.
Jag trodde att Tom skulle få panik.
Jag trodde att Tom skulle gripas av panik.
Jag trodde att Tom skulle råka i panik.
Jag trodde att Tom skulle bli panikslagen.
Jag trodde aldrig att Tom skulle sluta prata.
Jag trodde aldrig att Tom skulle hålla käften.
Snälla rätta mig när jag gör fel.
Fastän de ser ut som det är Carlos och Juan inte enäggstvillingar, bara bröder.
Jag vill inte översätta den här meningen.
Jag vill inte översätta denna mening.
Du är det vackraste flickan jag någonsin sett.
Hon är lång och smal.
Han reste under antaget namn.
Han reste under fingerat namn.
Han reste under täcknamn.
Fortsätt arbeta.
Du kan inte backa ur.
Du får inte backa ur.
Du kan inte hoppa av.
Du får inte hoppa av.
Du får inte smita.
Tom kan inte sitta i bilen längre än tio minuter innan han blir åksjuk.
Vi kan inte dödas.
Vi får inte dödas.
Tom kan inte lämnas ensam.
Jag kan inte förstå att jag precis sköt mig själv.
Jag kan inte fatta att vi äntligen klarade det.
Du kan inte skylla på mig.
Du får inte skylla på mig.
Jag kan inte bryta mig loss.
Jag kan inte bryta mig fri.
Jag kan inte knäcka den här koden.
Jag kan inte röra det ur fläcken.
Jag kan inte flytta på det.
Man kan inte köpa respekt.
Du kan inte köpa respekt.
Du får inte ringa Tom.
Jag kan inte sjunga en ren ton.
Jag kan inte ändra på det.
Du kan inte ändra på Tom.
Ni kan inte ändra på Tom.
Man kan inte ändra på Tom.
Jag kan inte ändra på vem jag är.
Jag kan inte komma just nu.
Jag kan inte komma i kväll.
Tom kan inte komma.
Jag kan inte delta.
Jag kan inte tävla.
Jag kan inte ställa upp.
Jag kan inte bekräfta det.
Jag kan inte bekräfta det.
Jag kan inte kontakta Tom.
Jag får inte kontakt med Tom.
Jag kan inte få kontakt med Tom.
Du kan inte kontrollera mig.
Ni kan inte kontrollera mig.
Man kan inte kontrollera mig.
Jag kan inte kontrollera Tom.
Jag kan inte övertyga Tom.
Jag kan inte heller dansa.
Jag kan inte dansa heller.
Jag kan inte dansa.
Jag kan inte hantera det här.
Du kan inte neka det.
Jag kan inte förneka det.
Tom kan inte göra någonting utan Marys hjälp.
Vi kan inte göra det nu.
Vi får inte göra det nu.
Jag kan inte göra det just nu.
Jag kan inte göra det i dag.
Jag klarar det inte i dag.
Vi kan inte göra det.
Jag kan inte göra det längre.
Jag kan inte göra det där heller.
Jag kan inte göra det nu.
Jag klara det inte nu.
Så kan Tom inte göra.
Tom kan inte göra så.
Tom kan inte göra det.
Tom får inte göra det.
Vi kan inte misslyckas.
Jag kan inte låtsas.
Jag kan inte bluffa det.
Jag kan inte fejka det.
Vi kan inte ge upp utan en kamp.
Du kan inte gå ut dit.
Du får inte gå ut dit.
Jag kan inte gå till polisen.
Du får inte skada Tom.
Du kan inte skada Tom.
Ni får inte skada Tom.
Ni kan inte skada Tom.
Jag kan inte bara stanna här.
Jag har ingen vodka.
Hon spelar Monopol.
Någon måste vara här för barnen.
Sikta. Skjut!
Fråga Tom.
Sluta!
Lägg av!
Var still.
Stilla.
Kom igen.
Kör vidare.
Ducka.
Fortsätt in.
Blidka mig.
Gör mig till viljes.
Låt det vara.
Låt den vara.
Lämna mig.
Lämna oss.
Gift dig med mig.
Stanna där du är!
Stanna där ni är!
Använd den här.
Använd det här.
Använd denna.
Använd detta.
Varna Tom.
Titta på hur jag gör det.
Titta hur jag gör det.
Kolla hur jag gör det.
Titta på mig.
Se på mig.
Titta på oss.
Se på oss.
Skriv till mig.
Du kan inte lämna mig.
Du får inte lämna mig.
Ni kan inte lämna mig.
Ni får inte lämna mig.
Jag kan inte lämna dig.
Vi kan inte låta Tom dö.
Jag kan inte låta dig göra det.
Jag kan inte låta er göra det.
Jag kan inte titta på Tom.
Du kan inte få oss att sluta.
Man kan inte stoppa tillbaka tandkräm i tuben.
Du kan inte sluta nu.
Du får inte sluta nu.
Ni får inte sluta nu.
Ni kan inte sluta nu.
Jag kan inte riktigt göra det.
Jag kan inte riktigt minnas.
Tom kan inte vägra.
Tom kan inte neka.
Tom kan inte säga nej.
Jag kan inte komma på texten.
Tom minns inte var.
Tom kan inte sjunga höga A.
Tom kan inte sjunga ett högt A.
Jag tål inte golf.
Jag står inte ut med sjukhus.
Jag klarar inte av lögnare.
Jag står inte ut med lögnare.
Tom kan inte stå still.
Jag klarar inte av att se blod.
Jag klarar inte av synen av blod.
Jag står inte ut med tanken på att förlora Tom som vän.
Jag står inte ut med tanken på att förlora dig för evigt.
Jag klarar inte av sådana här filmer.
Jag klarar inte av sådan här musik.
Jag kan inte riskera någonting.
Jag kan inte ta några risker.
Vi kan inte prata nu.
Du kan inte lita på någon.
Vi kysstes bara.
Jag vet bara vad Tom berättade för mig.
Jag ville bara prata med Tom.
Jag väger bara 45 kilo.
Jag var bara där en gång.
Jag gick bara dit en gång.
Jag önskar bara att jag kunde vara så lycklig som du verkar.
Jag önskar bara att jag kunde hjälpa er alla.
Om det bara var så enkelt.
Jag önskar bara att det var så enkelt.
Om det bara vore så enkelt.
Jag önskar bara hjälpa.
Jag vill bara vara till hjälp.
Jag önskar bara att Tom vore här.
Jag önskar bara att Tom kunde vara här.
Vad vill du ska hända?
Vad vill du berätta för oss?
Vad vill du titta på?
Var är resten av pengarna?
Vad hände med resten av maten?
Du ljuger!
Vi kan inte bevisa att Tom ljuger, men vi är ganska säkra på att han gör det.
Tom ljuger. Jag gjorde inte det som han sa att jag gjorde.
Det är tydligt att någon ljuger.
Jag undrar vem av er som ljuger.
Tom ligger på en stor sten.
Tom ligger på backen.
Tom ligger i sängen.
Tom ligger på rygg.
Offret låg med ansiktet ned i mattan.
Du berättar inte sanningen.
Vart går du oftast och klipper dig?
Hon har köpt en ny dator.
Regnet stod som spön i backen.
Jag har tappat bort min penna.
Jag ser fram emot sommarlovet.
Tom spelar på hästar.
Tom kunde inte tro på det som hänt.
Tom tog tag i Marys hand.
Tom skadade knät.
Du kommer inte kunna övertala Tom att göra det där.
Jag tänkte på Tom.
Jag trodde att jag hörde musik.
Jag trodde att jag hörde dig.
Jag trodde att jag kände dig.
Jag trodde att jag såg ett spöke.
Jag trodde att jag sa åt dig att inte komma.
Jag tyckte jag sa åt dig att inte stå i vägen för mig.
Jag trodde att jag förstod dig.
Jag trodde att jag var ensam.
Jag trodde att jag var trevlig.
Jag trodde att jag var lyckligt.
Jag tyckte att jag var lycklig.
Jag trodde att jag var i tid.
Jag trodde att jag förlorat dig,
Jag trodde att jag förlorat er.
Jag trodde att det var ett skämt.
Jag tänkte att det var värt ett försök.
Jag trodde att det skulle vara värt det.
Jag tänkte att det skulle vara värt det.
Jag trodde att fienden hade dödat Tom.
Jag trodde att Tom erkände.
Jag trodde att Tom hade stuckit.
Jag trodde Tom vad en fullständig idiot.
Jag trodde att Tom var död.
Jag trodde Tom var död.
Jag trodde att vi kunde prata.
Jag trodde att vi var bästa vänner.
Jag trodde att du hade en överenskommelse med Tom.
Jag trodde att du hatade Tom.
Jag trodde att du gillade mig.
Jag trodde du gillade mig.
Jag trodde att ni gillade mig.
Jag trodde ni gillade mig.
Jag trodde att du tyckte om mig.
Jag trodde du tyckte om mig.
Jag trodde att ni tyckte om mig.
Jag trodde ni tyckte om mig.
Jag trodde att du gillade Tom.
Jag trodde att du tyckte om Tom.
Jag trodde att ni två var lika gamla.
Jag trodde att du åkte hem.
Jag trodde att du gick hem.
Jag trodde att ni åkte hem.
Jag trodde att ni gick hem.
Jag trodde att du var Tom.
Jag trodde att du skulle hålla med.
Jag trodde att du åkt.
Jag trodde att du skulle gilla det.
Jag trodde att du skulle gilla den.
Jag trodde att du skulle tycka om det.
Jag trodde att du skulle tycka om den.
Jag trodde att ni skulle gilla den.
Jag trodde att ni skulle gilla det.
Jag trodde att ni skulle tycka om den.
Jag trodde att ni skulle tycka om det.
New York är en av de största städerna i världen.
Tom verkar vara en idiot.
Sjön ser ut som ett hav.
De skyndade sig ut ur rummet.
Det gick ju smärtfritt.
Han drar ifrån.
Jag tror fortfarande på kärleken.
Hon stod käpprak.
Jag skulle vilja få ett allvarsord med dig.
Vi skattade oss lyckliga som överlevde.
När man talar om trollen!
När man talar om trollen så står de i farstun.
Det är inte lätt att lösa problemet.
Återvänd till skeppet.
Jag behöver de här pengarna.
Jag behöver dessa pengar.
Vilket skepp var du på?
Ombord på vilket skepp var du?
Var är skeppet nu?
Varför är du på det här skeppet?
Varför är ni på det här skeppet?
Varför är ni på detta skepp?
Varför är du på detta skepp?
Fienden förstörde många av våra skepp.
Jag rörde ingenting.
Varför tar du på min flickvän?
Varför rör du min flickvän?
Vi försökte att kontakta det andra skeppet.
Skulle du kunna vara tyst, tack?
Orkanen Sandy är på väg.
Han tog sin tid.
Deras skepp ligger fortfarande i hamn.
Vilket skepp kom Tom med?
Vilket skepp kommer du med?
Jag är kapten över detta skepp.
Jag undrar vem som namngav detta skepp.
Vi går tillbaka till skeppet.
Vi måste gå tillbaka till skeppet.
Vårt skepp blev inte skadat i striden.
Jag undrar vart det där skeppet är på väg.
Var kom det där skeppet ifrån?
Vi ses igen när vi är tillbaka på skeppet.
Skeppet börjar sakta att röra på sig.
Det här är en bild på skeppet som jag var på.
Tom berättade för oss att det var ett gammalt skepp.
Vi kommer att söka genom hela skeppet.
Vi ska söka genom hela skeppet.
Tom föddes på ett skepp.
Vem är kapten över det här skeppet?
Vem är kapten över detta skepp?
Skeppet har inte ens dockat än.
De såg antagligen vårt skepp komma in i hamnen.
Tom sa att han läste en bok om det här skeppet.
Jag minns att jag var på ett skepp när jag var bara fem år gammal.
Hur långt borta tror du att det där skeppet är?
Skeppet genomsöktes noggrant, men inga illegala droger hittades.
När ska skeppet anlända?
När ska skeppet komma fram?
Jag har rätt att vara på det här skeppet.
Skeppet var inte redo för strid.
Var är kaptenen för det här skeppet?
Varför är du inte redan ombord på skeppet?
Jag kände att jag bara var tvungen att komma av skeppet.
Du blev tillsagd att stanna på skeppet.
Det här är det bästa skepp som jag någonsin varit på.
Tom tittade ut genom fönstret på skeppet som kom in i hamnen.
Det är ingen på det här skeppet förutom oss.
Hur många människor var ombord på det där skeppet?
Är Tom fortfarande kapten över ditt skepp?
Vi blev tillsagda att stanna på skeppet.
Jag har precis kommit hem.
Jag har precis kommit hem.
Min far är på promenad i parken.
Hon säger att hon inte dejtar någon just nu, men jag tror inte på henne.
Tom dricker inte öl hemma.
Om en dörrvakt bär ditt bagage, glöm inte att ge honom dricks.
De simmade.
Vi drack en hel del.
Vi drack mycket.
Var är min tidning?
Låt inte den här informationen läcka ut.
Det jag skrev är inte engelska.
Om det inte låter engelskt är det inte engelska.
Känner du någon som var på det där skeppet som sjönk?
Tror du att vi borde överge skeppet?
Jag gillar manga.
Jag gillar serieböcker.
Jag gillar tecknat.
Kriget tog slut 1954.
Varför lär jag mig isländska?
Varför läser jag isländska?
Varför studerar jag isländska?
De vill att vi ska tro att vi lever i en demokrati.
Jag skickade ett brev till Steina på isländska.
Jag hittade en mycket intressant hemsida som lägger fram fullständiga texter om isländska sagor, av vilka några också är översatta till engelska och danska.
Confucius sade: "Den som inte dricker te är en dåre."
När jag fantaserade fram fantasibilder fantaserade jag att min fantasiförmåga fantaserade alla bilderna. Tänk dig att ens fantasiförmåga fantaserar fram fantasier som man inte ens kan fantasera om.
Han har möjligheten att arbeta!
Hon har möjligheten att arbeta!
Den här jakten är väldigt dyr.
Den här yachten är väldigt dyr.
Denna lustjakt är väldigt dyr.
Vad ska du göra på Halloween?
Är du redo för Halloween?
Är det något särskilt?
Är det något särskilt som du vill?
Är det något särskilt som du vill höra?
Är det något särskilt som du vill titta på?
Är det något särskilt som du vill ha att äta?
Är det något särskilt som du vill ha att dricka?
Jag arbetade ihjäl mig i det där projektet.
Jag vill egentligen bara skaffa vänner.
En bra mening är bättre än två dåliga.
Det där är faktiskt riktigt elakt.
Vi klagar alltid.
Hur ser du om någon är en löpare?
Hur vet du om någon är en löpare?
De är oss på spåren!
Det här är ganska exakt.
Rör er inte!
Tamy upptäckte ett misstag i meningsbyggnaden.
Jag fick min välförtjänta lön.
Middagen är klar!
Middagen är färdig!
Lunchen är klar!
Vart går han?
Hur var Hawaii?
Han vill ha en iPad.
Hon vill ha en fjärde generationens iPad.
Han gav sin karriär som poet ett brått slut.
Tigern rymde från djurparken.
En av tigrarna rymde från djurparken.
En av tigrarna rymde från zoot.
Hans fru är svenska.
Du borde läsa en sådan bok som han läser just nu.
Mina planer misslyckades rejält.
Mina planer misslyckades kapitalt.
Regeringens politik misslyckades kapitalt.
Alla har rätt till sin egen åsikt. Men ibland är det bättre att hålla den för sig själv.
Tom är en av mina vänner.
Tom är en av mina närmsta vänner.
Jag är Toms vän.
Jag saknar mina vänner.
Jag är Marys pojkvän.
Jag var tillsammans med vänner hela förra natten.
Jag har en flickvän.
Jag blev Toms vän.
Jag fick just en vän.
Jag kanske är din enda vän.
Jag önskar att jag hade fler vänner.
Jag har en vän vid namn Tom.
Jag har en vän vars namn är Tom.
Jag har en vän som heter Tom.
Jag sov inte bra i natt, så jag har inte så mycket energi i dag.
Vad skrattar du åt?
Jag vill bara vara din vän, ingenting mer.
Jag har inga nära vänner.
Jag har alla de vänner som jag behöver.
Jag värdesätter vår vänskap.
Jag har ingen flickvän.
Jag har bara femtio med rep.
Vad ska du göra på fredag?
Vad ska du göra under sommarlovet?
Vad ska du göra på sommarlovet?
Tom tar en snabb joggingtur runt kvarteret varje morgon innan frukost.
Fattigdom lär en att äta bröd utan smör.
Jag vill ha två korv med bröd med mycket peppar.
En infraröd stråle består av elektromagnetisk strålning.
Han fjällade en fisk.
Vad är skillnaden mellan amerikansk och brittisk engelska?
Ser du den mustaschprydda mannen där borta?
Det är ett väldigt farligt system.
Det måste finnas ett mönster.
Tom är en urusel dansare.
Se till att Tom ringer mig.
Hämta Tom.
Ta tag i den där.
Hugg tag i Tom.
Visa hur man gör det där.
Visa mig.
Jag kysste henne på pannan.
Det här är en snuskig film.
Är det här Paris eller Marseille?
Vänta. Skjut inte än.
Sluta skjuta!
Tom alltid på sig en hatt.
Tom har nästan alltid på sig en hatt.
Tom har ofta på sig en hatt.
Tom har ofta på sig en hatt.
Tom har ibland på sig en hatt.
Tom har sällan på sig hatt.
Tom bär sällan hatt.
Tom har sällan på sig hatt.
Tom bär sällan hatt.
Tom har nästan aldrig på sig hatt.
Tom bär nästan aldrig hatt.
Tom har inte alltid hatt på sig.
Tom bär inte alltid hatt.
Tom har inte ofta på sig hatt.
Tom bär inte ofta hatt.
Tom har vanligtvis inte på sig hatt.
Tom har på sig hatt nästan varje dag.
Tom har på sig hatt varje dag.
Tom har inte hatt på sig varje dag.
Jag glömde min egen födelsedag.
Faktiskt så hittade jag på det där.
Faktiskt så är jag inte särskilt säker.
Kan du tro att detta faktiskt händer?
Hände det verkligen?
Sa verkligen Tom det?
Trodde du verkligen det?
Gav du verkligen Tom pengar?
Läste du verkligen det?
Såg du verkligen Tom?
Jag jobbar faktiskt här.
Jag gick faktiskt aldrig på högskola.
Jag såg det faktiskt inte själv.
Jag trodde inte att Tom faktiskt skulle prova det.
Jag har faktiskt aldrig träffat Tom.
Jag såg det faktiskt aldrig.
Jag är faktiskt en väldigt bra förare.
Jag är faktiskt ganska seriös.
Jag har faktiskt kul ikväll.
Jag är faktiskt ganska trött.
Jag är faktiskt väldigt upptagen.
Jag är faktiskt väldigt lycklig.
Jag är faktiskt här för att hjälpa dig.
Jag har faktiskt aldrig varit full.
Jag har faktiskt aldrig spelat golf.
Händer detta verkligen?
Det är faktiskt inte riktigt så enkelt.
Det var faktiskt inte så illa.
Det låter som om du faktiskt menar det.
Det var faktiskt mitt fel.
Det är faktiskt mycket enklare än vad det ser ut.
Det är faktiskt en bra poäng.
Det är faktiskt inte sant.
Det är faktiskt ganska smart.
Det är faktiskt bra nyheter.
Det är därför jag är här, faktiskt.
Tom trodde faktiskt på dig.
Tom gjorde faktiskt det han sa att han skulle göra.
Tom kom faktiskt på det själv.
Tom fick faktiskt Mary till att dansa med honom.
Tom gillar faktiskt Mary.
Tom spelar faktiskt inte mycket.
Tom pratar faktiskt inte mycket Franska.
Tom är faktiskt väldigt bra på att laga mat.
Tom var faktiskt inte där.
Toms party var ganska roligt, faktiskt.
Vi behöver faktiskt inte göra det nu.
Vem var det som faktiskt genomförde operationen?
Jag har inga böcker att läsa.
Jag har ingenting att läsa.
Jag har inget att skriva med.
Jag har ingenstans att gå.
Jag har inga kläder att använda.
Jag har inga rena kläder att använda.
Snälla gå ut härifrån genast.
Snälla gå ut ur mitt kontor genast.
Jag kan inte låta dem fånga mig.
Jag kan inte låta dem fånga dig.
Han sov i bilen.
Jag behöver förstå vad denna mening betyder.
Jag har bott här hela mitt liv.
Kan jag få tala med henne?
Vi gick ut på en promenad efter frukost.
Han är inte alltid glad.
Öppna inte lådan än.
Öppna inte presenten än.
Jag tror inte att kärlek finns.
Jag kan inte ens göra en omelett.
Jag kan inte förstå någonting av det han säger.
Han gick upp tidigt för att han skulle komma i tid till tåget.
Jag är din bror.
Jag är er bror.
Du ska alltid skydda dina ögon från direkt solljus.
Att bli klar med detta jobbet innan tisdag kommer att vara enkelt.
Att blir klar med det här jobbet innan tisdag kommer att bli enkelt.
Att bli klar med det här jobbet innan tisdag kommer att vara enkelt.
Att bli klar med detta jobb innan tisdag kommer att bli enkelt.
Att bli klar med detta jobb innan tisdag kommer att vara enkelt.
Han gillar grönsaker, framförallt vitkål.
Det vore bättre om du inte åt innan du gick till sängs.
Kan du snälla säga hur lång du är och din vikt?
Kan du snälla säga hur lång du är och hur mycket du väger?
Snälla ge mig ett plåster och lite medicin.
Jag mår inte bra. Snälla ge mig lite medicin.
Min far har slutat röka på grund av sin hälsa.
Min far har slutat röka för sin hälsas skull.
Tack för att du accepterade min vänförfrågan på Facebook.
Och det här är min sida.
Och detta är min sida.
Hon kunde inte sluta le.
Tom sa alltid att han ville lära sig spela mahjong.
Toms mamma sa alltid till honom att han borde äta mer grönsaker.
Du kanske har rätt.
Det var väldigt roligt.
Det var riktigt roligt.
Det var hemskt roligt.
Det var extremt roligt.
Det var ganska roligt.
Det var nästan roligt.
Det var inte roligt alls.
Klockan är nästan sju. Vi måste gå till skolan.
Min engelsklärare rekommenderade mig att läsa dessa böcker.
Min engelsklärare rekommenderade mig att läsa de här böckerna.
Jag har fyra datorer, men två av dem är så gamla att jag inte använder dem längre.
Regler är regler.
Hon är så jävla charmig!
Hur var din dag idag?
Släpp ankaret!
Ju mer pengar vi har, desto mer vill vi ha.
Jag tvättade min T-shirt.
Hur träffade du din partner?
Jag sovde väldigt bra.
Mitt te är för sött.
Tom spenderade hela dagen med att designa en hemsida åt en ny kund.
Tom brukade röka två paket cigaretter varje dag.
Toms fru gillar inte när han röker i vardagsrummet.
Jag skrattade väldigt mycket när jag såg det där.
Jag skyller på ditt skägg.
Vill du ha te eller något?
Har du blivit en ängel?
Är han inte söt när han är arg?
Jag svär att jag aldrig ska göra det igen.
Ärligt talat, jag är inte särskilt imponerad av hans idée.
Dimman var så tjock att jag inte kunde se vart jag var påväg.
Jag är förföljd.
Jag ska lära ut Esperanto i mitt land.
John tände en tändsticka.
Du glömde att dividera med X här.
Vad gjorde han efter det?
Vänta en sekund. Detta telefonsamtalet kan vara viktigt.
Röstade du?
Vem blir den nästa presidenten av USA?
Vem röstade du på?
Vem kommer att vinna i Ohio?
Folk ändras. Det finns inte mycket du kan göra åt det.
Jag vet precis vem Tom tänker gifta sig med.
Jag tror att hon är ärlig
Jag tror hon är ärlig.
Jag tror han är ärlig.
Läs inte vad som är i brevet. Bara ge det till Tom.
Jag matade hunden.
Min hund bet Tom.
Detta är väldigt lätt.
Jag hoppas att något bra händer innan dagen är över.
Jag är riktigt trött. Idag gick jag alldeles för mycket.
Har du dina biljetter?
Jag har en hund som kan springa snabbt.
Detta är total demagogi.
Alla dörrar i huset var stängda.
Ingen står över lagen.
Ställ inga frågor.
Vad gjorde du i skolan idag?
Vem åt den sista kakan?
Det är hemligt.
Har du lärt dig din läxa?
Fråga inte, bara gör det.
Jag ställde inga frågor.
Jag ville bara ställa en fråga.
Låt mig fråga en fråga.
Snälla fråga inte en sådan fråga.
När jag läste till jurist sa mina lärare åt mig att aldrig ställa en fråga som jag inte visste svaret på.
När jag läste till advokat sa mina lärare åt mig att aldrig ställa en fråga som jag inte visste svaret på.
Skulle du ha något emot att jag ställer en fråga?
Du frågar ofta frågor som jag inte kan svara på.
Gillar du sött te?
Vad för fråga är det där?
Njuter du av det här?
Njuter du av detta?
Njuter ni av det här?
Njuter ni av detta?
Är du road av det här?
Är du road av detta?
Är ni roade av det här?
Är ni roade av detta?
Tyckte du om det där?
Njöt du av det där?
Tyckte du om matchen?
Hade du roligt på matchen?
Tyckte du om föreställningen?
Hade du roligt på föreställningen?
Tyckte du om rundturen?
Hade du kul på turnén?
Tyckte du om rundvandringen?
Njuter du av att förlora?
Hon är ganska söt.
Han pratade aldrig om det.
Hon pratade aldrig om det.
Han vill inte prata om det.
Jag kommer att behöva din hjälp.
Kan du japanska?
Kan ni tala japanska?
Jag har inte tid att läsa böcker.
Han har aldrig varit i Amerika.
Du ser precis ut som din pappa.
Snälla lämna.
Jag förstår.
Min far är stolt över det faktum att han aldrig varit i en trafikolycka.
Varför är tjejer så komplicerade?
Tjejer är inte komplicerade. Män är simpla.
Jag antar att vi har gjort ett helt okej jobb eftersom ingen har klagat.
Problemet med den svenska animationsbranschen är att den i stort sett är icke-existerande.
Själv föredrar jag vodka, men jag har inget emot att ta en likör ibland.
Min flickvän är helt tokig i Forever 21, men det är åtminstone billigt.
Varje gång jag sätter på mikrovågsugnen så slutar mitt Wi-Fi att fungera, det är extremt irriterande.
Jag skulle vilja ha ett ord med dig.
Jag är riktigt stolt över dig.
En god mandellikör skulle allt sitta bra nu.
Hellre död än röd.
Hellre död än röd.
Kan jag räkna med dig?
Kan jag lita på dig?
Mobbning är så klart ett allvarligt problem, men samtidigt måste vi inse att en nollvision här är omöjlig.
Det ska du ha jävligt klart för dig!
Visst, min mamma är prostituerad, men på den ljusa sidan så har vi åtminstone någonstans att bo.
Robotarna kommer att ta över en dag, det kan du vara säker på.
Visst älskar jag Finland, men jag står inte ut med finnarna.
Du kanske inte tittar så mycket på TV?
Din mamma är en riktig snuskhummer, Pelle. Jag orkar inte med hennes insinuationer!
Bra jobbat, gubbar.
Vill du att jag ska ringa polisen?
Min man blev så ställd att han tappade sina bilnycklar.
Jag har inte mycket till övers för Hollywoods superhjältefilmer.
Driver du med mig?
Du måste skämta!
Jag håller inte med, det är inte rasistiskt att använda ordet "ras".
Det finns ju vissa uttryck som numera bara används ironiskt.
Ingen har bett dig att hålla med, men du kan väl åtminstone acceptera att det finns personer som har andra åsikter än dig?
Fet chans.
Jaha, det var ju just en stor överraskning också.
Nä, säger du det?
Visst kan det vara traumatiskt, men än sen?
Jag litar inte på politiker.
Båda mina föräldrar var arbetslösa, men det hindrade dem inte från att ta väl hand om mig och mina 23 syskon.
Snubben som står i hörnet där borta kan röka upp en cigarett på mindre än en minut.
På 80-talet var det minsann andra bullar som gällde.
Jag tar en kebabpizza special, med blandad sås.
Svårt att tro, men så är det.
Du måste skämta!
Är jag i trubbel?
Han bad om ett glas vatten.
Tom är död.
Tom är rädd.
Tom är en hippie.
Tom är ursinnig.
Tom är gift.
Tom saknas.
Tom arbetar.
I sina böcker rasade han ofta mot regeringen och dess politik.
Vi kan inte göra det.
Vem dog?
Vem har dött?
Hans kropp hittades aldrig.
Tom beslutade sig för att börja med flugfiske.
Ett sätt att minska antalet fel i Tatoebas korpus skulle vara att uppmuntra människor att endast översätta till sina modersmål.
Den här boken är unik på många sätt.
Jag läste ett brev.
Jag läser ett brev.
Jag vill vinna.
Jag vill ha en öl.
Vi vill rösta.
Ingen vill ha ett krig.
Jag vill bara veta.
Jag vill inte leka.
Jag vill inte spela.
Jag vill inte vila.
Jag vill inte ha dig här.
Jag vill inte ha er här.
Jag vill bara hjälpa er.
Jag vill bara hjälpa dig.
Jag vill ha ett par handskar.
Jag vill ha en förklaring.
Jag vill ha tillbaka mina tjugo dollar.
Jag vill att du kommer tillbaka till Boston.
Jag vill inte störa Tom.
Jag vill bara vara med dig.
Berätta för Tom vad du vill göra.
Tom ville inte tala med mig.
Tom ville inte prata med mig.
Tom sa att han ville vara här.
Tom sade att han ville vara här.
Du vill ha dom här grejerna, inte sant?
Vill du gå någon annanstans?
Jag vill inte att någon ska bli skadad.
Jag vill inte gå till jobbet idag.
Jag vill inte höra några ursäkter.
Tom vill inte prata med dig.
Varför skulle någon vilja göra det?
Jag vill inte göra några misstag.
Jag ville att Tom skulle känna sig som hemma.
Hördu, jag vill inte förlora mitt jobb.
Ingen av oss vill gifta sig.
Jag var nära att dö av en hjärtattack.
Vill du att jag ska hålla ett öga på Tom åt dig?
Jag vill att du kommer tillbaka nästa vecka.
Om du inte vill att jag ska åka, så gör jag det inte.
Hon är en drama queen.
Ungarna spelar Duck Hunt.
Barnen spelar Duck Hunt.
Det kan vi inte göra.
Flodens övre lopp är mycket vackert.
Ljuger du för mig?
Jag bor på Malta.
Jag vill ha en förklaring och jag vill ha den nu!
Jag vill ha svar och jag vill ha dem nu!
Tom är skadad.
Kineserna vet inte att jag inte är mänsklig.
Du förtjänar mer.
Jag vill verkligen inte lämna barnen ensamma nu.
Jag vill att du går på mötet imorgon.
Han tittade på en svensk film.
Jag tittade på en svensk film i går kväll.
Greta Garbo var en svensk skådespelare.
Kameran som du köpte är bättre än min.
Det sägs att han är den bästa tennisspelaren.
Jag vill inte att det ska finnas några lögner mellan oss.
Om du vill köpa ett koppel, gå till en zooaffär.
Om du tänker döda mig så vill jag veta varför.
Jag vill veta vad som är roligt.
Jag vill veta vad som är så roligt.
Jag vill veta vad det är som är roligt.
Jag vill veta vad det är som är så roligt.
Varför skulle Tom vilja hjälpa oss?
Till följd av konstant hunger och utmattning dog hunden till slut.
Jag vill veta exakt vad det är som händer.
Jag vet att du inte ville att Tom skulle åka in i fängelse.
Jag bestämde mig för att jag inte ville ha mer med Tom att göra.
Jag ser inget problem med detta.
Han kan tala franska och engelska.
Hon säljer en ny hatt.
Vi pratade om diverse olika ämne.
Jag vill bara kunna besöka mina barn när jag så önskar.
Jag vill bara kunna besöka mina barn när jag vill.
Om du vill prata, prata.
Om du vill prata så prata.
Om du vill prata, prata då.
Jag skulle vilja gå och sova nu.
Jag var så lycklig på den tiden.
Det var nästan som en dröm.
Jag hoppas att det här är början på en vacker vänskap.
Det låter som om du är upptagen.
Tom har svimmat.
Du måste inte bestämma dig just nu.
Du borde vara försiktigare nästa gång.
Du borde vara noggrannare nästa gång.
Ni borde vara försiktigare nästa gång.
Ni borde vara noggrannare nästa gång.
Allt måste handskas med väldigt försiktigt.
Jag tycker att du är lite för försiktig.
Jag tror att du är lite för försiktig.
Jag tycker att du är lite för noggrann.
Jag tror att du är lite för noggrann.
Tom är här.
Det där var riktigt kul. Gör det igen!
Det där var riktigt roligt. Gör det igen!
Vi klarar oss.
Var snäll och spika igen fönstren.
Läs detta först.
Läs det här först.
Det var fortfarande riktigt varmt, trots att solen hade sjunkit ganska lågt.
Mark tog sina saker och gick.
Tycker du att jag är larvig?
Tycker ni att jag är larvig?
Jag planerar att tala fler än 20 språk år 2015.
Huset tillhör honom.
Ingen kommer att klandra dig.
Ingen kommer att beskylla dig.
Ingen kommer att klandra er.
Ingen kommer att beskylla er.
Något fruktansvärt har hänt.
Någonting fruktansvärt har hänt.
Är det något fel på dina ögon?
Jag tror att vi glömde någonting.
Har du ingenting att göra?
Har inte du något att göra?
Har ni ingenting att göra?
Har inte ni något att göra?
Å, det är en världslig sak!
Du måste kämpa mot den tendensen hos dig.
När blir det klart?
Tom går till skolan till fots.
Vi är från Ryssland.
Vad är den turkiska motsvarigheten till meditation?
Han var tvungen att lämna skolan för att han var fattig.
Kasta inte bort den här tidningen!
Han ringde mig.
Vi upptäckte en hemlig passage.
Vem?
Jag tror inte att de kommer att acceptera dessa villkor.
Mannen som ringde för en timme sedan var Frank.
I byn finns inga tjuvar.
Jag visste inte att hon har ett barn.
Det är kallt ute.
Ingen skall överleva.
Ingen kommer att överleva.
Ingen får gå dit.
Var är min son?
Jag nyser hela tiden.
Tom älskar Mary.
Jag älskar min stad.
Välkommen, John! Vi väntade på dig.
Och vad sade de till mig?
Och vad sa de till mig?
Och vad berättade de för mig?
Vänligen, mata inte djuren!
Skriv aldrig orden "borsjtj" och "sjtji" på tyska!
Jag förstår att Volapük är ett bra språk.
Berings sund avskiljer Asien från Nordamerika.
Inte här!
Tom är adopterad.
Tom är alert.
Tom är på alerten.
Tom är uppmärksam.
Tom är snabb i vändningarna.
Tom är vid liv.
Tom är ensam.
Tom är allena.
Tom är för sig själv.
Tom är road.
Tom är arg.
Tom är ängslig.
Tom har anlänt.
Tom är vaken.
Tom blöder.
Tom bluffar.
Tom är uttråkad.
Tom är genialisk.
Tom fuskar.
Tom är gladlynt.
Tom är glad av sig.
Tom är munter.
Tom håller på att kvävas.
Tom är bekymrad.
Tom har erkänt.
Tom är förvirrad.
Tom är vid medvetande.
Tom är vid sans.
Tom är övertygad.
Tom lagar mat.
Tom har rätt.
Tom är tokig.
Tom är galen.
Tom gråter.
Tom är farlig.
Tom är döv.
Tom har dött.
Tom är annorlunda.
Tom är skild.
Tom är i våningen under.
Tom är i nedre våningen.
Tom drömmer.
Tom drunknar.
Tom är full.
Tom dör.
Tom är tidig.
Tom äter.
Tom är förlovad.
Tom har rymt.
Tom är känd.
Tom är snabb.
Tom är tjock.
Tom är fet.
Tom är orädd.
Tom är oförskräckt.
Tom är smutsig.
Tom är lortig.
Tom är färdig.
Tom är stollig.
Tom är hispig.
Tom är knäpp.
Tom är fri.
Tom är vänlig.
Tom är rolig.
Tom är glad.
Tom är borta.
Tom har åkt.
Tom har gått.
Tom är snål.
Tom sörjer.
Tom är ostadig på benen.
Tom är groggy.
Tom är skyldig.
Tom är oförarglig.
Tom är ofarlig.
Tom är halsstarrig.
Tom är hårdnackad.
Tom är egensinnig.
Tom är styvsint.
Tom hjälper till.
Tom hjälper.
Tom är hemma.
Tom är hemlös.
Tom har hemlängtan.
Tom är hungrig.
Tom är imponerad.
Tom är mentalsjuk.
Tom är sinnessjuk.
Tom är vansinnig.
Tom är vanvettig.
Tom skämtar.
Tom skrattar.
Tom har åkt.
Tom haltar.
Tom är ensam.
Tom har tur.
Tom är lyckligt lottad.
Tom ljuger.
Tom är arg.
Tom är elak.
Tom packar.
Tom målar.
Tom är artig.
Tom är framfusig.
Tom är framåt.
Tom har sagt upp sig.
Tom vilar.
Tom är pensionerad.
Tom har kommit tillbaka.
Tom har rätt.
Tom är ledsen.
Tom är säker.
Tom är blyg.
Tom är sjuk.
Tom är tyst.
Tom är ärlig.
Tom är smart.
Tom är hög.
Tom är konstig.
Tom är sträng.
Tom är stark.
Tom är trött.
Tom är uppe.
Tom väntar.
Tom är svag.
Tom vinner.
Tom är orolig.
Tom är ängslig.
Tom är bekymrad.
Tom har fel.
Tom är ung.
Vi förlorade.
Vi lovade.
Vi överlevde.
Vi väntade.
Vi kommer att överleva.
Vi ska vinna.
Vi kommer att vinna.
Han sköt först!
Hennes hobby är bodybuilding.
Tom kör.
De kommer att attackera.
De kommer att anfalla.
Det är utpressning.
Ta min.
Ta mitt.
Tag min.
Tag mitt.
Jag är ursinnig.
Jag är rasande.
Jag är skild.
Jag ser.
Klä på dig.
Klä på er.
Hitta Tom.
Vänta inte.
Stanna inte.
Stirra inte.
Stå inte.
Tala inte.
Prata inte.
Le inte.
Sjung inte.
Skrik inte.
Spring inte!
Rör dig inte!
Titta inte.
Ljug inte.
Hoppa inte!
Slåss inte.
Fuska inte.
Öl är gott.
Var tolerant.
Var toleranta.
Var hänsynslös.
Var hänsynslösa.
Tom är stark.
Jag valde mellan två alternativ.
Ibland är det försent att be om ursäkt.
Var god och tag plats!
Det är alltid värt ett försök.
Kyrkan står mitt i byn.
Jag vet knappt någonting alls.
Strävan efter sanning är beundransvärd.
Att sträva efter sanning är beundransvärt.
Ge aldrig upp!
Han är ett matvrak.
Hon är en storätare.
Hon är ett matvrak.
Regimen störtades till slut.
Jag gör mitt bästa.
Förresten såg jag honom igår.
Typisk tjejsnack!
Var snäll och avbryt mig inte.
Tack för ditt mejl!
Det vore kul att träffas snart igen.
Livet kunde vara en dröm.
Livet skulle kunna vara en dröm.
Djur kan inte särskilja mellan sant och falskt.
Låt oss vara ärliga!
Allting var förberett långt i förväg.
Du är annorlunda.
Den är tom.
Det är tomt.
Jag hittade min borttappade plånbok.
Vi får inte många besökare här nere.
Jag vet att jag är "osvensk". Och det tänker jag fortsätta att vara. Lagom är inte bäst; bäst är bäst!
Hur många äpplen då?
Han är dum som ett spån.
En skola i Storbritannien har frångått läroböcker till förmån för iPads i klassrummet.
Kinesiska tidningar övervakas av regeringen som behåller rätten att ändra innehåll för att passa den rådande partilinjen.
Brott lönar sig inte i längden.
Kriminalitet lönar sig inte i längden.
Kriminalitet lönar sig inte i det långa loppet.
Kriminalitet lönar sig inte på lång sikt.
Hon har något emot rödhåriga.
Talar ni bulgariska?
Talar ni bulgariska?
Denna förordning träder i kraft från och med nästa år.
Du gissade rätt. Boken var fortfarande i bilen.
Mitt löfte att komma nästa måndag håller fortfarande.
Han läser en bok.
Jag ser ut som en ren.
Körsbären blomstrar i april.
Han kommer snart.
Där är en pojke.
Klandra inte mig! Jag har inte något att göra med den där videon.
Skyll inte på mig. Jag har ingenting att göra med den där videon.
Det är svårt att tala offentligt.
Jag är fri som en fågel.
Jag ångrar att jag inte åkte dit.
Jag ångrar att jag inte gick dit.
Var bor du just nu?
Var bor ni just nu?
Den här motorn ger ibland upp andan.
Klockan var fem i ett när jag gick till sängs.
Klockan var fem i ett när jag gick och la mig.
Klockan var fem i ett när jag gick och lade mig.
Hon var fem i ett när jag gick till sängs.
Hon var fem i ett när jag gick och la mig.
Hon var fem i ett när jag gick och lade mig.
Var nu inte så skadeglad!
Låt inte folk göra dig galen över pengar, hår och kläder.
Skulle du vilja ha ett glas vatten?
Är din fru kvar i Amerika?
Är din fru fortfarande i Amerika?
Du var min räddare i nöden.
Vi hörs.
Ursäkta, var ligger posten?
Ni vet att vi inte har så mycket tid just nu.
Jag tror att den här killen menar allvar.
Men det är ju absurt.
Han har gått ur tiden.
Jag har inte ätit soppan och jag kommer inte att göra det.
Han är absolutist.
Detta är inte acceptabelt.
Vilken är din favoritactionrulle?
Det var en av mitt livs mest makalösa upplevelser.
Min far, farfar, farfars far och farfars farfar hade alla samma namn som jag.
Hon är aggressiv.
Om du tror att det var mitt fel är du inne på fel spår.
Erfarenheten räknas.
Det är likartat.
Det är liknande.
Det är likt.
Den är liknande.
Den är lik.
Vid midnatt skall jag gå fram genom Egypten, och allt förstfött i Egyptens land skall dö.
Jag vet att det inte är lätt.
Han är mycket oförskämd.
Han är väldigt oförskämd.
Vilken underbar trädgård!
Kosta vad det kosta vill.
Vill du ha en snigel på ögat?
Damaskus ligger i Syrien.
Det går upp för mig.
Inga skämt, tack!
Sköt om dig!
Hon tittade på några klänningar och valde ut den dyraste.
Boken är på bordet.
Sluta prata om min familj.
Försökt inte att fly från ansvar.
Sådant händer.
Koncentrera dig på ditt uppdrag!
Koncentrera dig på vårt uppdrag!
Det knackar på dörren.
Boken kostar fyra dollar.
Jag gick upp för en timme sen.
Varför har koalor ingen navel?
Vem är allsångsledare i år?
Han går som en anka.
Jag är utledsen på det.
Jag är urless på det.
Jag är utled på det.
Om det blir några svårigheter, ring mig!
Tom hade en benägenhet att titta bort när han blev tilltalad.
Dessa tvillingbröder är lika som bär.
Vad tänker du på just nu?
De har inga barn, så vitt jag vet.
Den här föreningen grundades för etthundraelva år sedan.
Egentligen ville vi gå på bio i lördags, men vi ångrade oss och stannade hemma.
När fadern kom hem, tittade jag på tv.
Här anrikar man malm.
Varför är du så arrogant?
Jag växte upp i en fattig familj.
Han kände medlidande med oss.
Jag är inte en pappersmugg.
Om det regnar i morgon, stannar vi hemma.
Var kan vi prata ostört?
Vad kan man göra åt det?
Jag är helt förvirrad.
Han har hår på bröstet.
Han har köpt ett bananfodral.
Det svider.
Hur många armar har en bläckfisk?
Hur många armar har en bläckfisk?
Vem äger dessa renar?
Jag vill inte prata om det just nu.
Krig är helvetet.
Var parkerade du bilen?
Jag glömde boken hemma.
Som pensionär är jag nu min egen chef - äntligen.
Hon tror att hon vet bäst.
Var inte så nyfikna!
Du är orättvis.
Ni är orättvisa.
Jag är upprörd.
Tom ringde.
Jag vinner.
Han är nykterist.
Jag är en sjusovare.
Jag är Döden.
Jag är här som turist.
Varför slutar du inte?
Varför slutar ni inte?
Hon har platinablont hår.
Äpplena är inte plockmogna än.
Han är en mycket attraktiv man.
Det beror på stolens storlek.
Det kan inte undvikas.
Vad tittar du på mig för?
Vad tittar ni på mig för?
Ni är alla bjudna.
Du ljuger ju bara.
Ni ljuger ju bara.
Du är bara nervös.
Du behövs inte.
Ni behövs inte.
Du är överflödig.
Du har rätt, Tom.
Du är Toms favorit.
Du måste arbeta snabbt.
Ni måste arbeta snabbt.
Det finns många arter av fiskmås som varierar i storlek.
Försök att inte äta för mycket.
Självklart tycker jag om det.
Gör inte om det.
Jag är egyptier.
Jag stod en stund och tittade på avgasröret.
Vi stötte på dem vid bussterminalen.
Tom tog någonting.
Vi ursäktar avbrottet.
Jag åkte aldrig fast.
Det visade sig att han visste allt om mig.
Tom och Mary har en mack ihop.
Jag köpte mackan på macken.
Tomten är inte till salu.
Tomten är inte till salu.
Det här trädet är inte ens i närheten av att vara det högsta i socknen.
Tom åkte tillbaka.
Tom gick tillbaka.
Tom försvann.
Vi har inget behov av assistans.
Vi är båda galna.
Vi är ganska säkra.
De köpte det.
De köpte den.
Flickan stirrade på dockan.
De ser förvirrade ut.
De ser bra ut.
De såg förskräckta ut.
De älskade det.
De älskade den.
De tog i hand.
De skakade hand.
De började dansa.
De började skjuta.
De började skjuta.
De gick ut.
De litar på dig.
De vill ha mig.
De ville ha bevis.
De blev tokiga.
De var falska.
Dom var utmärkta.
De var hjältar.
De var mina.
De blev mördade.
De mördades.
De var perfekta.
Skyskrapan förväntas sjunka ner i myren.
Varför tror du att jag tänker på dig?
Det är bara en teori.
De ville inte lyssna.
Sover du?
Är vi inte vänner?
Ring mig senare.
Ring polisen.
Ring snuten.
Vann du?
Vann ni?
Var inte barnslig.
Jag gick inte.
Jag stjäl inte.
Jag känner mig sårbar.
Jag fastnade.
Jag tappade kontrollen.
Jag behövde det här.
Jag behövde dig.
Jag behövde er.
Är han död?
Fetma är en nationell epidemi.
Jag arbetade.
Jag flyttar inte.
Jag flyttar mig inte.
Jag flyttar inte på mig.
Jag kommer att följa dig.
Är allt där?
Smittar det?
Det kommer aldrig att hända.
När du är i Rom, bete dig som romarna.
Det är inte billigt.
Det där är inte billigt.
Vilken lättnad!
Vilken relief!
Vem hatar dig?
Vilka är det som hatar dig?
Vem hatar er?
Vilka är det som hatar er?
Du kan inte se.
Du får inte se.
Du förtjänar det här.
Du verkar förvånad.
Ni verkar förvånade.
Äh, tyst med dig.
Hon grät sig till sömns.
Din katt är tjock.
Er katt är tjock.
Jag kan inte använda vänster hand på grund av gipset.
Ge mig något att skriva på.
Ge mig något att signera.
Jag håller med Tom.
Hur träffade du honom?
Han går vanligtvis hem klockan fem.
Vi har inget annat val.
Elefanter är majestätiska djur.
Det är den bästa vi har.
Ibland är det viktigt att fatta ett beslut snabbt.
Nu eller aldrig.
Det skulle vara trevligt om jag kunde resa till Japan.
Hörde du mig inte?
Hörde ni mig inte?
Vi väntade på båten i många timmar.
Vi åker om en vecka idag.
Du ser ut som en liten flicka i den klänningen.
Kvinnan är rik, men mannen är fattig.
Jag dricker inte champagne.
Jag ska inte förråda Tom.
Jag kommer inte att behöva dig.
Jag kommer inte att behöva er.
Äta bör man, annars dör man. Äta gör man, ändå dör man.
Ingenting är sant; allt är tillåtet.
Tom bröt mot reglerna.
Tom är min brorson.
Tom är min systerson.
Du har stavat mitt namn fel.
Ni har stavat mitt namn fel.
Du har felstavat mitt namn.
Ni har felstavat mitt namn.
Du har stavat fel på mitt namn.
Ni har stavat fel på mitt namn.
Titta inte på kameran.
Jag vet inte riktigt än.
Ett slukhål har bildats mitt i motorvägen.
Det är där jag kommer att vara.
Jag kan inte läsa skrivstil, så kan du vara snäll och texta?
En katt låg och sov i bastrumman.
Åt du frukost?
Åt ni frukost?
Du är en idiot!
Han har ett stort ego.
Vem förrådde oss?
Han kör utan körkort.
Jag kan göra det härifrån.
Jag kan inte låta det hända.
Var inte en sådan surpuppa!
Jag kunde inte fortsätta ljuga för Tom.
Jag kunde inte stoppa Tom.
Vi blev goda vänner.
Vi drack lite vin.
Han lärde sig att skriva siffror innan han kom till skolan.
Jag tappade kontrollen.
Och vad gör vi nu?
Hon har självmordstankar.
Jag köpte en ny handväska.
Hjälp mig bygga färdigt den här sorkstegen så ska jag bjuda dig på middag.
Jag går till skolan på lördag.
Han var synligt nervös.
Jag var tvungen att hämta någonting från mitt rum.
Han är en sefardisk jude.
Detta är min dator.
Håll tummarna för mig!
Du är så ondskefull!
Ni är så ondskefulla!
Du har blivit tjock.
Jag har många samtal att ringa.
Jag har många beslut att fatta.
Jag har inte sovit något vidare.
Jag har bra dagar och dåliga dagar.
Jag har aldrig röstat.
Jag vet inte om vi kan hjälpa dig eller inte.
Jag kan inte minnas att jag har bett om din hjälp.
Jag kommer inte att följa med dig.
Jag tänker inte lyssna på dig.
Jag är nykter.
Använd en skalpell, inte en yxa.
Jag ska vila mig lite.
Tack! Du är fantastisk!
Tack! Ni är fantastiska!
Skynda dig, tåget stannar bara här en kort stund.
Skynda er, tåget stannar bara här en kort stund.
Har du något käk?
Jag vet att du är arg.
Du håller på att bli lat!
Ni håller på att bli lata!
Jag lät mina känslor fördunkla mitt omdöme.
Jag ljög för dig.
Jag ljög för er.
Han är inte arg.
Han är inte galen.
Varför är hunden här?
Jag förlorade allt som jag hade.
Jag har gjort kaffe åt dig.
Jag gjorde kaffe åt dig.
Jag har gjort kaffe åt er.
Jag gjorde kaffe åt er.
Jag fick dig att känna dig obekväm, inte sant?
Jag fick dig att skratta, eller hur?
Jag fick er att skratta, eller hur?
Jag gör dig nervös, inte sant?
Jag gör er nervösa, inte sant?
Jag behöver en bil.
Jag låtsades arbeta.
Jag hoppas verkligen att du har rätt.
Jag hoppas verkligen att ni har rätt.
Jag minns allt du säger till mig.
Kan du tala esperanto?
Kan ni tala esperanto?
Hur fattar du dina beslut?
Hur fattar ni era beslut?
Jag sa att det var ok.
Jag såg Tom för mindre än en timme sen.
Jag såg Tom för mindre än en timme sedan.
Jag tror att Tom och John är enäggstvillingar.
Jag tycker att vi borde vänta.
Hon är gift med en tandläkare.
Han är gift med en tandläkare.
Har du ätit frukost?
Har ni ätit frukost?
Mannen åt bröd.
Har du ätit frukost?
Jag vill inte att arbeta under dessa betingelser.
Han begick många synder i sin ungdom.
Om jag då hade kunnat tala franska, hade jag inte fått några problem.
Talar Tom flytande franska?
Ursäkta mig, jag har en förfrågan.
Jag var där ensam i början, men sedan kom Liisa och Liisas nya vän.
Det var trevligt att göra ingenting.
Liisa är en aktiv och energisk ung kvinna.
Använd ditt självförtroende, men aldrig visa upp den för mycket!
Det internationella språket interlingue offentliggjordes 1922 under namnet Occidental.
Tre av mina barn dog.
Tror du att det kommer att regna idag?
Tror ni att det kommer att regna idag?
Du har helt rätt.
Ni har helt rätt.
Jag låtsades arbeta.
Vad sägs om en promenad på stranden?
Smör görs av mjölk.
Det finns en annan möjlighet också.
Du är avskedad!
Var ligger hotellet?
Betty dödade sin egen mor.
Jag tror att jag har gjort mitt; det är din tur nu.
Skällde hunden?
Hunden har hållit på och skälla.
Kan jag kyssa dig?
Får jag kyssa dig?
Din fråga är ologisk.
Skratta inte!
Liisa hade inte en aning om vad hon skulle göra.
Låt mig ge dig ett råd.
Det är inte blod. Det är tomatsås.
Markku satte sitt liv på spel för att rädda Liisa.
Och återigen var han hur full som helst.
Har du någonsin sett Buckingham Palace?
Välkommen till Wikipedia, den fria encyklopedin som alla kan redigera.
Varför kan Tom inte komma?
Hon pratar inte bara flytande engelska utan också flytande franska.
Varning! Vått golv.
Är detta en hingst eller ett sto?
Jag var inte medveten om att Tom hade gjort det.
Jag är i princip lika kvalificerad som Tom.
Tom tände bordslampan.
Jag ska aldrig glömma Toms ansikte.
Jag ska berätta sanningen.
Tom kunde inte öppna dörren.
Tom moppar golvet.
Jag får inte gå härifrån.
Jag går till kyrkan.
Min kniv är vass.
Det är ingen hemlighet.
Jag tänker, alltså är jag.
Jag vill inte se dum ut.
Jag vill inte verka dum.
Jag var lärare.
Det var aldrig svårt för oss att hitta något att prata om.
Varför har du inte klänning på dig?
Ta på dig en klänning då.
Alkohol löser inga problem.
Vad undersöker en sovjetolog?
Vad studerar en sovjetolog?
Livet är som en stor huvudväg.
Kvinnan äter bröd.
Det här bordet är vitt.
Jag kommer från Turkiet.
Det ligger en apelsin på bordet.
Jag är rädd för höjder.
Jag är höjdrädd.
Det finns ett fel i meningen.
Abonnenten du försöker nå kan inte ta ditt samtal just nu. Vänligen försök igen senare.
Åt du något?
Jag brände pappret.
Jag brände papperet.
Ingången till toaletten är mycket smutsig.
Hur många gånger måste jag säga det till dig?
Jag är inte läkare.
Kärleken är en viktig sak.
Europa är en kontinent.
Mitt hjärta blöder.
Jag skall gå till stranden.
Jag ska gå till stranden.
Det där är ett hjärta.
Jag skall äta äpplet.
Jag gick inte till skolan.
Jag skall gå till parken.
Jag ska gå till parken.
Jag har blå ögon.
Jag har röda ögon.
Talar du arabiska?
Hassan gick till skolan.
Han är min dubbelgångare.
Vill du ha fisk?
Jag talar arabiska.
Katten är under bordet.
Han återvänder till sitt hem.
Han åt äpplet.
Jag har ett hjärta.
Jag har en katt.
Jag skall läsa boken.
Jag ska läsa boken.
Jag är studerande.
Vetenskapen är viktig för våra liv.
Jag tror inte att två språk är tillräckligt.
Tom släckte lampan på nattduksbordet.
Tom och Mary var dom två sista att ge sig av.
Tom och Mary var på Johns begravning.
Tom arbetade deltid.
Tom ser verkligen ledsen ut.
Varför är dom rädda?
Var är dina barn?
Var är era barn?
Vi hade våra skäl.
Vad är vi skyldiga?
Det är ovanligt.
Jag lokaliserar programvaran.
Jag kan inte äta.
Jag kan äta.
Jag kan leva utan vatten.
Det nya huset ligger här.
Det här är mitt hus.
Du sover i mitt rum.
Jag frågar henne en fråga.
Emily frågade en fråga.
Jag återvände från skolan.
Det finns en katt i lådan.
Jag öppnar en låda.
Han kan simma.
Hon kan simma.
Jag köpte henne en vacker klänning.
Jag drack kaffet.
Emily kan simma.
Det här är en hönsfågel.
Min penna är i min hand.
Ditt blod är rött.
Jag går och lägger mig klockan tio.
Jag bor i Qatar.
Jag går till jobbet klockan sju.
Jag går och lägger mig klockan tio.
Jag skrev inte ett brev.
Jag drack inte vattnet.
Hur länge tänker du stanna här i Brasilien?
Emily skriver ett brev.
Te är en populär dryck över hela världen.
Jag kan inte förstå.
Du kommer att förstå att jag berättar sanningen.
Jag sjunger en sång.
Jag sjunger en skön sång.
Bilen är blå.
Jag måste göra min läxa.
Du måste göra din läxa.
Jag äter en bok.
Vi vann tävlingen!
Jag förstår dina ord.
Har du en ordbok?
Jag behöver en bättre ordbok.
Jag vill lära mig svenska.
Jag återvände till huset.
Det här äpplet är rödare.
Vad är din blodgrupp?
Stockholm är Sveriges huvudstad.
Sveriges huvudstad är Stockholm.
Katten sover på bordet.
Vilken skola är bäst?
Jag gick till sjukhuset.
Alla rören frös förra vintern.
För ögonblicket har vi större problem.
Just nu, har vi större problem.
Brevet är skrivet av flickan.
Någon stal mitt körkort.
Jag delar inte din åsikt.
Jag hörde åskdundret, men såg inte blixten.
Låt oss spatsera litet på stranden.
Detta fält är inte väl odlat.
Älskar du henne?
Jag har lärt mig något från den här boken.
Hon hade gått till skolan.
Staden ligger vid havsstranden.
Jag kan älska det.
Vi behöver köpa vinäger.
Hon öppnade dörren.
Jag talar tyska.
Frukosten serveras klockan sju.
Grattis!
Jag funderade på planen.
Räven byter pälsen men inte lasterna.
Ett fruktansvärt kaos härskar i vardagsrummet.
Hon slöt sina ögon.
Han är elva år gammal.
Fången befanns skyldig.
Jag har ett dåligt samvete.
Bar båda hjälmar?
Rökning är förbjudet.
Den här filmen är ett mästerverk.
Han är sällan hemma.
Han bodde i Azerbajdzjan i 4 år.
Då ska jag se vad jag kan göra!
Påven Francis återvänder till Rio år 2016.
Om ni sticker oss, blöda vi icke?
Om jag bara hade bett om ditt råd.
Toms far är en berömd konstnär.
Han kommer att vara ledig imorgon.
Jag förmodar att han kommer.
Jag skulle vilja ha en gaffel.
Jag skulle vilja skicka ett rekommenderat brev.
Hon ville avsäga sig sitt amerikanska medborgarskap.
Jag har många språkböcker.
Jag vill vara ett barn.
Jag vill inte leva med dig.
Den här byggnaden ska byggas i staden.
Jag talar lite franska.
Har ni sett den här?
Vampyren suger mitt blod.
Hon ljög.
Alla djur är lika.
Jag har en vit katt.
Heather tror mig.
Jag spelar i trädgården.
Det är inte möjligt.
Jag vill gifta mig med Heather.
Jag talar om ditt handlande.
Jag talar om ditt agerande.
Vem sitter vanligtvis på åsnebänken?
Vem sitter vanligtvis på åsnebänken?
Vem sitter vanligtvis på åsnebänken?
Det är förnedrande för henne.
Afrika är mänsklighetens vagga.
Hur många delfiner finns det på detta oceanarium?
Hon hatade vanilj.
Jag måste vara försiktig.
Snälla sluta!
Emily är en gottegris.
Jag ska berätta det för Emily.
Emily ska berätta det för Melanie.
Jag kramade Emily.
Emily kramade mig.
Min engelska är inte god.
Min engelska är inte bra.
Jag vill tala engelska.
Det är felaktigt.
Emily vill arbeta i ett stort företag.
Jag skulle vilja köpa en hund.
Det finns en pojke i det här rummet.
Det finns en hund i det här rummet.
Du kan inte ersätta kommat med en punkt i den här meningen.
Jag ser fram emot det.
Du sa till honom.
Vi säljer skor.
Han varnade dig.
Hon varnade dig.
Hur kan speglar vara sanna om våra ögon inte är äkta?
Hon kopierade en mening.
Jag läser den här tidningen.
Hon förklarade ett skämt.
Hon översatte en dikt.
Hon tvättade en matta.
Hon vattnade ett träd.
Hon vann en telefon.
Hon bar en mask.
Hon skrev en kort berättelse.
Emily skrev meningen.
Jag åkte till Norge.
Jag åkte till Sverige.
Jag åkte till Danmark.
Vi gick till stranden.
Hon sjöng en sång.
Du borde gå till en läkare.
Är du inte riktigt klok?
På golvet stod två par skor.
Du har fått det du ville, lämna mig ifred nu.
Hon försöker begå självmord.
Varför i helvete lever du såhär, Tom?
Jag dricker vatten i köket.
Jag har frågor.
Hon kan spela gitarr.
Är du rädd för höjder?
Jag måste lära mig ett språk.
Behöver du något?
Behöver ni någonting?
Jag behöver en bok att läsa.
Han kan ruttna i helvetet.
Jag vill skriva en bok.
Tom har en ko.
Emet gillar inte den kvinnan.
Markku verkade glatt överraskad.
Vi vill att regeringen ska tjäna hela befolkningen.
Emet ogillar den där kvinnan.
Sjärnorna ser mycket vackra ut i kväll.
Vi har ingen dotter.
Tänker du ligga i sängen hela dagen, eller?
Jag läser inte så många böcker som jag gjorde tidigare.
Fanns inga moln på himlen.
Blomman är röd.
Han lagade en middag för henne.
Vi hjälpte dem.
Jag lovar att säga till om jag ser något passande.
Solenergitekniken är kostnadseffektiv nuförtiden.
Jag måste åka till Danmark i morgon.
Jag är i Ryssland.
