ställ konen på den röda cirkeln på cirkeln 
ta konen på cirkeln 
ta blocket
ta ett block 
ställ en röd kon på cirkeln 
ställ blocket på den blåa cirkeln på cirkeln 
ställ den blåa konen på den blåa cirkeln 
ställ den blåa konen på den röda cirkeln 
ställ det blåa blocket på den röda cirkeln 
ställ det röda blocket på den röda cirkeln 
ställ den röda konen på den blåa cirkeln på cirkeln 
ta den blåa konen på den röda cirkeln 
ta den blåa konen på den blåa cirkeln 
ställ blocket på cirkeln på den röda cirkeln 
ta konen 
ta blocket 
ställ blocket på cirkeln på cirkeln 
ta det blåa blocket  
ta ett blått block 
ta konen på den röda cirkeln 
ställ blocket på den röda cirkeln 
ställ blocket på cirkeln på den röda cirkeln 
ta konen 
ställ den röda konen på cirkeln 
ställ konen på cirkeln på den röda cirkeln 
ställ det blåa blocket på den blåa cirkeln 
ta blocket på cirkeln 
ta det röda blocket 
ta den röda konen på cirkeln 
ställ konen på den röda cirkeln på den röda cirkeln 
ställ blocket på den röda cirkeln 
ta det blåa blocket 
ställ blocket på den röda cirkeln 
ställ den blåa konen på den röda cirkeln 
ställ det blåa blocket på den blåa cirkeln 
ta konen 
ställ konen på den röda cirkeln på cirkeln 
ta det blåa blocket 
ställ konen på cirkeln på den röda cirkeln 
ställ konen på cirkeln på cirkeln 
ta blocket på den röda cirkeln 
ta blocket 
ställ den röda konen på den röda cirkeln 
ta det blåa blocket 
ta blocket 
ta det blåa blocket 
ställ den blåa konen på cirkeln 
ställ blocket på cirkeln på den blåa cirkeln 
ställ konen på den röda cirkeln på den röda cirkeln 
ta det röda blocket 
ställ den blåa konen på den blåa cirkeln 
ställ det röda blocket på den blåa cirkeln 
ställ konen på cirkeln 
ställ den blåa konen på cirkeln på cirkeln 
ställ konen på den röda cirkeln på cirkeln 
ställ det blåa blocket på den röda cirkeln 
ställ konen på den röda cirkeln på cirkeln 
ta konen 
ställ den blåa konen på cirkeln 
ta konen 
ställ den blåa konen på den röda cirkeln på cirkeln 
ställ den röda konen på den röda cirkeln 
ställ blocket på den blåa cirkeln 
ta konen på cirkeln 
ställ konen på cirkeln på cirkeln 
ställ blocket på den röda cirkeln 
ta blocket på cirkeln 
ställ det blåa blocket på den blåa cirkeln 
ta det röda blocket 
ta konen 
ställ konen på cirkeln 
ta den röda konen 
ställ konen på cirkeln på den röda cirkeln 
ställ den röda konen på cirkeln 
ställ konen på cirkeln på den röda cirkeln 
ta det röda blocket på den blåa cirkeln 
ta det röda blocket 
ta blocket 
ställ det röda blocket på den blåa cirkeln 
ställ blocket på cirkeln på cirkeln 
ställ konen på cirkeln på den röda cirkeln 
ställ det röda blocket på cirkeln 
ställ konen på cirkeln 
ställ blocket på den blåa cirkeln på cirkeln 
ställ konen på den röda cirkeln 
ta det röda blocket 
ställ det röda blocket på cirkeln på den blåa cirkeln 
ställ konen på den röda cirkeln på cirkeln 
ställ den blåa konen på den blåa cirkeln 
ställ blocket på cirkeln 
ställ konen på cirkeln 
ta det blåa blocket 
ställ den röda konen på cirkeln på cirkeln 
ställ blocket på den röda cirkeln 
ställ den blåa konen på den röda cirkeln 
ställ den röda konen på cirkeln 
ställ den blåa konen på den röda cirkeln på cirkeln 
ta den blåa konen 
ställ det röda blocket på den blåa cirkeln 
ställ det blåa blocket på den röda cirkeln 
ställ konen på den blåa cirkeln 
ta det blåa blocket 
ställ en pil på den röda cirkeln på cirkeln
ta pilen på cirkeln
ta ett block
jag ställer en röd kon på cirkeln
hon ställer en röd kon på cirkeln
jag ställer mitt block på den blåa cirkeln på cirkeln
hon ställer en blå pil på den blåa cirkeln
han ställer sin blåa pil på den röda cirkeln
han ställer ett blått block på den röda cirkeln
hon ställer sitt röda blocket på den röda cirkeln
ställ den röda konen på den blåa cirkeln på cirkeln
ta den blåa konen på den röda cirkeln
ta en blå kon på den blåa cirkeln
han ställer sitt block på cirkeln på den röda cirkeln
han tar konen
jag tar blocket
jag ställer mitt block på cirkeln på cirkeln
jag tar det blåa blocket
ta konen på den röda cirkeln
jag ställer blocket på hennes röda cirkeln
jag ställer blocket på hans cirkel på hennes röda cirkel
hon tar sin kon
jag ställer den röda pilen på min cirkel
ställ konen på cirkeln på den röda cirkeln
ställ det blåa blocket på den blåa cirkeln
ta blocket på cirkeln
ta det röda blocket
ta den röda konen på cirkeln
ställ en pil på den röda cirkeln på den röda cirkeln
ställ blocket på en röd cirkel
ta det blåa blocket
ställ blocket på den röda cirkeln
ställ den blåa konen på den röda cirkeln
ställ det blåa blocket på den blåa cirkeln
ta konen
ställ pilen på den röda cirkeln på cirkeln
ta det blåa blocket
ställ pilen på cirkeln på den röda cirkeln
ställ konen på cirkeln på cirkeln
ta blocket på den röda cirkeln
ta ett block
ställ den röda konen på den röda cirkeln
ta det blåa blocket
ta blocket
ta det blåa blocket
ställ den blåa konen på cirkeln
ställ blocket på cirkeln på den blåa cirkeln
ställ konen på den röda cirkeln på den röda cirkeln
ta det röda blocket
ställ en blå kon på en blå cirkel
ställ ett rött block på en blå cirkel
ställ konen på en cirkel
ställ den blåa konen på cirkeln på cirkeln
ställ en pil på den röda cirkeln på cirkeln
ställ ett blått block på den röda cirkeln
ställ konen på den röda cirkeln på cirkeln
ta konen
ställ en blå pil på cirkeln
ta en kon
ställ en blå pil på den röda cirkeln på en cirkel
ställ den röda konen på den röda cirkeln
ställ blocket på den blåa cirkeln
ta konen på cirkeln
ställ konen på cirkeln på cirkeln
ställ blocket på den röda cirkeln
ta blocket på cirkeln
ställ det blåa blocket på den blåa cirkeln
ta det röda blocket
ta pilen på cirkeln
ställ konen på cirkeln
ta en röd pil
ställ den röda pilen på cirkeln
ställ pilen på cirkeln på den röda cirkeln
ställ pilen på cirkeln på den röda cirkeln
ställ den blåa pilen på den blåa cirkeln
ställ den röda pilen på cirkeln på cirkeln
ställ en pil på den röda cirkeln
ställ den röda konen på en cirkel
ta en pil
